magic
tech sky130A
magscale 1 2
timestamp 1640630825
<< obsli1 >>
rect 1104 493 583803 701777
<< obsm1 >>
rect 566 8 583815 701808
<< metal2 >>
rect 8114 703200 8170 704000
rect 24306 703200 24362 704000
rect 40498 703200 40554 704000
rect 56782 703200 56838 704000
rect 72974 703200 73030 704000
rect 89166 703200 89222 704000
rect 105450 703200 105506 704000
rect 121642 703200 121698 704000
rect 137834 703200 137890 704000
rect 154118 703200 154174 704000
rect 170310 703200 170366 704000
rect 186502 703200 186558 704000
rect 202786 703200 202842 704000
rect 218978 703200 219034 704000
rect 235170 703200 235226 704000
rect 251454 703200 251510 704000
rect 267646 703200 267702 704000
rect 283838 703200 283894 704000
rect 300122 703200 300178 704000
rect 316314 703200 316370 704000
rect 332506 703200 332562 704000
rect 348790 703200 348846 704000
rect 364982 703200 365038 704000
rect 381174 703200 381230 704000
rect 397458 703200 397514 704000
rect 413650 703200 413706 704000
rect 429842 703200 429898 704000
rect 446126 703200 446182 704000
rect 462318 703200 462374 704000
rect 478510 703200 478566 704000
rect 494794 703200 494850 704000
rect 510986 703200 511042 704000
rect 527178 703200 527234 704000
rect 543462 703200 543518 704000
rect 559654 703200 559710 704000
rect 575846 703200 575902 704000
rect 570 0 626 800
rect 1674 0 1730 800
rect 2870 0 2926 800
rect 4066 0 4122 800
rect 5262 0 5318 800
rect 6458 0 6514 800
rect 7654 0 7710 800
rect 8758 0 8814 800
rect 9954 0 10010 800
rect 11150 0 11206 800
rect 12346 0 12402 800
rect 13542 0 13598 800
rect 14738 0 14794 800
rect 15934 0 15990 800
rect 17038 0 17094 800
rect 18234 0 18290 800
rect 19430 0 19486 800
rect 20626 0 20682 800
rect 21822 0 21878 800
rect 23018 0 23074 800
rect 24214 0 24270 800
rect 25318 0 25374 800
rect 26514 0 26570 800
rect 27710 0 27766 800
rect 28906 0 28962 800
rect 30102 0 30158 800
rect 31298 0 31354 800
rect 32402 0 32458 800
rect 33598 0 33654 800
rect 34794 0 34850 800
rect 35990 0 36046 800
rect 37186 0 37242 800
rect 38382 0 38438 800
rect 39578 0 39634 800
rect 40682 0 40738 800
rect 41878 0 41934 800
rect 43074 0 43130 800
rect 44270 0 44326 800
rect 45466 0 45522 800
rect 46662 0 46718 800
rect 47858 0 47914 800
rect 48962 0 49018 800
rect 50158 0 50214 800
rect 51354 0 51410 800
rect 52550 0 52606 800
rect 53746 0 53802 800
rect 54942 0 54998 800
rect 56046 0 56102 800
rect 57242 0 57298 800
rect 58438 0 58494 800
rect 59634 0 59690 800
rect 60830 0 60886 800
rect 62026 0 62082 800
rect 63222 0 63278 800
rect 64326 0 64382 800
rect 65522 0 65578 800
rect 66718 0 66774 800
rect 67914 0 67970 800
rect 69110 0 69166 800
rect 70306 0 70362 800
rect 71502 0 71558 800
rect 72606 0 72662 800
rect 73802 0 73858 800
rect 74998 0 75054 800
rect 76194 0 76250 800
rect 77390 0 77446 800
rect 78586 0 78642 800
rect 79690 0 79746 800
rect 80886 0 80942 800
rect 82082 0 82138 800
rect 83278 0 83334 800
rect 84474 0 84530 800
rect 85670 0 85726 800
rect 86866 0 86922 800
rect 87970 0 88026 800
rect 89166 0 89222 800
rect 90362 0 90418 800
rect 91558 0 91614 800
rect 92754 0 92810 800
rect 93950 0 94006 800
rect 95146 0 95202 800
rect 96250 0 96306 800
rect 97446 0 97502 800
rect 98642 0 98698 800
rect 99838 0 99894 800
rect 101034 0 101090 800
rect 102230 0 102286 800
rect 103334 0 103390 800
rect 104530 0 104586 800
rect 105726 0 105782 800
rect 106922 0 106978 800
rect 108118 0 108174 800
rect 109314 0 109370 800
rect 110510 0 110566 800
rect 111614 0 111670 800
rect 112810 0 112866 800
rect 114006 0 114062 800
rect 115202 0 115258 800
rect 116398 0 116454 800
rect 117594 0 117650 800
rect 118790 0 118846 800
rect 119894 0 119950 800
rect 121090 0 121146 800
rect 122286 0 122342 800
rect 123482 0 123538 800
rect 124678 0 124734 800
rect 125874 0 125930 800
rect 126978 0 127034 800
rect 128174 0 128230 800
rect 129370 0 129426 800
rect 130566 0 130622 800
rect 131762 0 131818 800
rect 132958 0 133014 800
rect 134154 0 134210 800
rect 135258 0 135314 800
rect 136454 0 136510 800
rect 137650 0 137706 800
rect 138846 0 138902 800
rect 140042 0 140098 800
rect 141238 0 141294 800
rect 142434 0 142490 800
rect 143538 0 143594 800
rect 144734 0 144790 800
rect 145930 0 145986 800
rect 147126 0 147182 800
rect 148322 0 148378 800
rect 149518 0 149574 800
rect 150622 0 150678 800
rect 151818 0 151874 800
rect 153014 0 153070 800
rect 154210 0 154266 800
rect 155406 0 155462 800
rect 156602 0 156658 800
rect 157798 0 157854 800
rect 158902 0 158958 800
rect 160098 0 160154 800
rect 161294 0 161350 800
rect 162490 0 162546 800
rect 163686 0 163742 800
rect 164882 0 164938 800
rect 166078 0 166134 800
rect 167182 0 167238 800
rect 168378 0 168434 800
rect 169574 0 169630 800
rect 170770 0 170826 800
rect 171966 0 172022 800
rect 173162 0 173218 800
rect 174266 0 174322 800
rect 175462 0 175518 800
rect 176658 0 176714 800
rect 177854 0 177910 800
rect 179050 0 179106 800
rect 180246 0 180302 800
rect 181442 0 181498 800
rect 182546 0 182602 800
rect 183742 0 183798 800
rect 184938 0 184994 800
rect 186134 0 186190 800
rect 187330 0 187386 800
rect 188526 0 188582 800
rect 189722 0 189778 800
rect 190826 0 190882 800
rect 192022 0 192078 800
rect 193218 0 193274 800
rect 194414 0 194470 800
rect 195610 0 195666 800
rect 196806 0 196862 800
rect 197910 0 197966 800
rect 199106 0 199162 800
rect 200302 0 200358 800
rect 201498 0 201554 800
rect 202694 0 202750 800
rect 203890 0 203946 800
rect 205086 0 205142 800
rect 206190 0 206246 800
rect 207386 0 207442 800
rect 208582 0 208638 800
rect 209778 0 209834 800
rect 210974 0 211030 800
rect 212170 0 212226 800
rect 213366 0 213422 800
rect 214470 0 214526 800
rect 215666 0 215722 800
rect 216862 0 216918 800
rect 218058 0 218114 800
rect 219254 0 219310 800
rect 220450 0 220506 800
rect 221554 0 221610 800
rect 222750 0 222806 800
rect 223946 0 224002 800
rect 225142 0 225198 800
rect 226338 0 226394 800
rect 227534 0 227590 800
rect 228730 0 228786 800
rect 229834 0 229890 800
rect 231030 0 231086 800
rect 232226 0 232282 800
rect 233422 0 233478 800
rect 234618 0 234674 800
rect 235814 0 235870 800
rect 237010 0 237066 800
rect 238114 0 238170 800
rect 239310 0 239366 800
rect 240506 0 240562 800
rect 241702 0 241758 800
rect 242898 0 242954 800
rect 244094 0 244150 800
rect 245198 0 245254 800
rect 246394 0 246450 800
rect 247590 0 247646 800
rect 248786 0 248842 800
rect 249982 0 250038 800
rect 251178 0 251234 800
rect 252374 0 252430 800
rect 253478 0 253534 800
rect 254674 0 254730 800
rect 255870 0 255926 800
rect 257066 0 257122 800
rect 258262 0 258318 800
rect 259458 0 259514 800
rect 260654 0 260710 800
rect 261758 0 261814 800
rect 262954 0 263010 800
rect 264150 0 264206 800
rect 265346 0 265402 800
rect 266542 0 266598 800
rect 267738 0 267794 800
rect 268842 0 268898 800
rect 270038 0 270094 800
rect 271234 0 271290 800
rect 272430 0 272486 800
rect 273626 0 273682 800
rect 274822 0 274878 800
rect 276018 0 276074 800
rect 277122 0 277178 800
rect 278318 0 278374 800
rect 279514 0 279570 800
rect 280710 0 280766 800
rect 281906 0 281962 800
rect 283102 0 283158 800
rect 284298 0 284354 800
rect 285402 0 285458 800
rect 286598 0 286654 800
rect 287794 0 287850 800
rect 288990 0 289046 800
rect 290186 0 290242 800
rect 291382 0 291438 800
rect 292578 0 292634 800
rect 293682 0 293738 800
rect 294878 0 294934 800
rect 296074 0 296130 800
rect 297270 0 297326 800
rect 298466 0 298522 800
rect 299662 0 299718 800
rect 300766 0 300822 800
rect 301962 0 302018 800
rect 303158 0 303214 800
rect 304354 0 304410 800
rect 305550 0 305606 800
rect 306746 0 306802 800
rect 307942 0 307998 800
rect 309046 0 309102 800
rect 310242 0 310298 800
rect 311438 0 311494 800
rect 312634 0 312690 800
rect 313830 0 313886 800
rect 315026 0 315082 800
rect 316222 0 316278 800
rect 317326 0 317382 800
rect 318522 0 318578 800
rect 319718 0 319774 800
rect 320914 0 320970 800
rect 322110 0 322166 800
rect 323306 0 323362 800
rect 324410 0 324466 800
rect 325606 0 325662 800
rect 326802 0 326858 800
rect 327998 0 328054 800
rect 329194 0 329250 800
rect 330390 0 330446 800
rect 331586 0 331642 800
rect 332690 0 332746 800
rect 333886 0 333942 800
rect 335082 0 335138 800
rect 336278 0 336334 800
rect 337474 0 337530 800
rect 338670 0 338726 800
rect 339866 0 339922 800
rect 340970 0 341026 800
rect 342166 0 342222 800
rect 343362 0 343418 800
rect 344558 0 344614 800
rect 345754 0 345810 800
rect 346950 0 347006 800
rect 348054 0 348110 800
rect 349250 0 349306 800
rect 350446 0 350502 800
rect 351642 0 351698 800
rect 352838 0 352894 800
rect 354034 0 354090 800
rect 355230 0 355286 800
rect 356334 0 356390 800
rect 357530 0 357586 800
rect 358726 0 358782 800
rect 359922 0 359978 800
rect 361118 0 361174 800
rect 362314 0 362370 800
rect 363510 0 363566 800
rect 364614 0 364670 800
rect 365810 0 365866 800
rect 367006 0 367062 800
rect 368202 0 368258 800
rect 369398 0 369454 800
rect 370594 0 370650 800
rect 371698 0 371754 800
rect 372894 0 372950 800
rect 374090 0 374146 800
rect 375286 0 375342 800
rect 376482 0 376538 800
rect 377678 0 377734 800
rect 378874 0 378930 800
rect 379978 0 380034 800
rect 381174 0 381230 800
rect 382370 0 382426 800
rect 383566 0 383622 800
rect 384762 0 384818 800
rect 385958 0 386014 800
rect 387154 0 387210 800
rect 388258 0 388314 800
rect 389454 0 389510 800
rect 390650 0 390706 800
rect 391846 0 391902 800
rect 393042 0 393098 800
rect 394238 0 394294 800
rect 395342 0 395398 800
rect 396538 0 396594 800
rect 397734 0 397790 800
rect 398930 0 398986 800
rect 400126 0 400182 800
rect 401322 0 401378 800
rect 402518 0 402574 800
rect 403622 0 403678 800
rect 404818 0 404874 800
rect 406014 0 406070 800
rect 407210 0 407266 800
rect 408406 0 408462 800
rect 409602 0 409658 800
rect 410798 0 410854 800
rect 411902 0 411958 800
rect 413098 0 413154 800
rect 414294 0 414350 800
rect 415490 0 415546 800
rect 416686 0 416742 800
rect 417882 0 417938 800
rect 418986 0 419042 800
rect 420182 0 420238 800
rect 421378 0 421434 800
rect 422574 0 422630 800
rect 423770 0 423826 800
rect 424966 0 425022 800
rect 426162 0 426218 800
rect 427266 0 427322 800
rect 428462 0 428518 800
rect 429658 0 429714 800
rect 430854 0 430910 800
rect 432050 0 432106 800
rect 433246 0 433302 800
rect 434442 0 434498 800
rect 435546 0 435602 800
rect 436742 0 436798 800
rect 437938 0 437994 800
rect 439134 0 439190 800
rect 440330 0 440386 800
rect 441526 0 441582 800
rect 442630 0 442686 800
rect 443826 0 443882 800
rect 445022 0 445078 800
rect 446218 0 446274 800
rect 447414 0 447470 800
rect 448610 0 448666 800
rect 449806 0 449862 800
rect 450910 0 450966 800
rect 452106 0 452162 800
rect 453302 0 453358 800
rect 454498 0 454554 800
rect 455694 0 455750 800
rect 456890 0 456946 800
rect 458086 0 458142 800
rect 459190 0 459246 800
rect 460386 0 460442 800
rect 461582 0 461638 800
rect 462778 0 462834 800
rect 463974 0 464030 800
rect 465170 0 465226 800
rect 466274 0 466330 800
rect 467470 0 467526 800
rect 468666 0 468722 800
rect 469862 0 469918 800
rect 471058 0 471114 800
rect 472254 0 472310 800
rect 473450 0 473506 800
rect 474554 0 474610 800
rect 475750 0 475806 800
rect 476946 0 477002 800
rect 478142 0 478198 800
rect 479338 0 479394 800
rect 480534 0 480590 800
rect 481730 0 481786 800
rect 482834 0 482890 800
rect 484030 0 484086 800
rect 485226 0 485282 800
rect 486422 0 486478 800
rect 487618 0 487674 800
rect 488814 0 488870 800
rect 489918 0 489974 800
rect 491114 0 491170 800
rect 492310 0 492366 800
rect 493506 0 493562 800
rect 494702 0 494758 800
rect 495898 0 495954 800
rect 497094 0 497150 800
rect 498198 0 498254 800
rect 499394 0 499450 800
rect 500590 0 500646 800
rect 501786 0 501842 800
rect 502982 0 503038 800
rect 504178 0 504234 800
rect 505374 0 505430 800
rect 506478 0 506534 800
rect 507674 0 507730 800
rect 508870 0 508926 800
rect 510066 0 510122 800
rect 511262 0 511318 800
rect 512458 0 512514 800
rect 513562 0 513618 800
rect 514758 0 514814 800
rect 515954 0 516010 800
rect 517150 0 517206 800
rect 518346 0 518402 800
rect 519542 0 519598 800
rect 520738 0 520794 800
rect 521842 0 521898 800
rect 523038 0 523094 800
rect 524234 0 524290 800
rect 525430 0 525486 800
rect 526626 0 526682 800
rect 527822 0 527878 800
rect 529018 0 529074 800
rect 530122 0 530178 800
rect 531318 0 531374 800
rect 532514 0 532570 800
rect 533710 0 533766 800
rect 534906 0 534962 800
rect 536102 0 536158 800
rect 537206 0 537262 800
rect 538402 0 538458 800
rect 539598 0 539654 800
rect 540794 0 540850 800
rect 541990 0 542046 800
rect 543186 0 543242 800
rect 544382 0 544438 800
rect 545486 0 545542 800
rect 546682 0 546738 800
rect 547878 0 547934 800
rect 549074 0 549130 800
rect 550270 0 550326 800
rect 551466 0 551522 800
rect 552662 0 552718 800
rect 553766 0 553822 800
rect 554962 0 555018 800
rect 556158 0 556214 800
rect 557354 0 557410 800
rect 558550 0 558606 800
rect 559746 0 559802 800
rect 560850 0 560906 800
rect 562046 0 562102 800
rect 563242 0 563298 800
rect 564438 0 564494 800
rect 565634 0 565690 800
rect 566830 0 566886 800
rect 568026 0 568082 800
rect 569130 0 569186 800
rect 570326 0 570382 800
rect 571522 0 571578 800
rect 572718 0 572774 800
rect 573914 0 573970 800
rect 575110 0 575166 800
rect 576306 0 576362 800
rect 577410 0 577466 800
rect 578606 0 578662 800
rect 579802 0 579858 800
rect 580998 0 581054 800
rect 582194 0 582250 800
rect 583390 0 583446 800
<< obsm2 >>
rect 572 703144 8058 703338
rect 8226 703144 24250 703338
rect 24418 703144 40442 703338
rect 40610 703144 56726 703338
rect 56894 703144 72918 703338
rect 73086 703144 89110 703338
rect 89278 703144 105394 703338
rect 105562 703144 121586 703338
rect 121754 703144 137778 703338
rect 137946 703144 154062 703338
rect 154230 703144 170254 703338
rect 170422 703144 186446 703338
rect 186614 703144 202730 703338
rect 202898 703144 218922 703338
rect 219090 703144 235114 703338
rect 235282 703144 251398 703338
rect 251566 703144 267590 703338
rect 267758 703144 283782 703338
rect 283950 703144 300066 703338
rect 300234 703144 316258 703338
rect 316426 703144 332450 703338
rect 332618 703144 348734 703338
rect 348902 703144 364926 703338
rect 365094 703144 381118 703338
rect 381286 703144 397402 703338
rect 397570 703144 413594 703338
rect 413762 703144 429786 703338
rect 429954 703144 446070 703338
rect 446238 703144 462262 703338
rect 462430 703144 478454 703338
rect 478622 703144 494738 703338
rect 494906 703144 510930 703338
rect 511098 703144 527122 703338
rect 527290 703144 543406 703338
rect 543574 703144 559598 703338
rect 559766 703144 575790 703338
rect 575958 703144 583444 703338
rect 572 856 583444 703144
rect 682 2 1618 856
rect 1786 2 2814 856
rect 2982 2 4010 856
rect 4178 2 5206 856
rect 5374 2 6402 856
rect 6570 2 7598 856
rect 7766 2 8702 856
rect 8870 2 9898 856
rect 10066 2 11094 856
rect 11262 2 12290 856
rect 12458 2 13486 856
rect 13654 2 14682 856
rect 14850 2 15878 856
rect 16046 2 16982 856
rect 17150 2 18178 856
rect 18346 2 19374 856
rect 19542 2 20570 856
rect 20738 2 21766 856
rect 21934 2 22962 856
rect 23130 2 24158 856
rect 24326 2 25262 856
rect 25430 2 26458 856
rect 26626 2 27654 856
rect 27822 2 28850 856
rect 29018 2 30046 856
rect 30214 2 31242 856
rect 31410 2 32346 856
rect 32514 2 33542 856
rect 33710 2 34738 856
rect 34906 2 35934 856
rect 36102 2 37130 856
rect 37298 2 38326 856
rect 38494 2 39522 856
rect 39690 2 40626 856
rect 40794 2 41822 856
rect 41990 2 43018 856
rect 43186 2 44214 856
rect 44382 2 45410 856
rect 45578 2 46606 856
rect 46774 2 47802 856
rect 47970 2 48906 856
rect 49074 2 50102 856
rect 50270 2 51298 856
rect 51466 2 52494 856
rect 52662 2 53690 856
rect 53858 2 54886 856
rect 55054 2 55990 856
rect 56158 2 57186 856
rect 57354 2 58382 856
rect 58550 2 59578 856
rect 59746 2 60774 856
rect 60942 2 61970 856
rect 62138 2 63166 856
rect 63334 2 64270 856
rect 64438 2 65466 856
rect 65634 2 66662 856
rect 66830 2 67858 856
rect 68026 2 69054 856
rect 69222 2 70250 856
rect 70418 2 71446 856
rect 71614 2 72550 856
rect 72718 2 73746 856
rect 73914 2 74942 856
rect 75110 2 76138 856
rect 76306 2 77334 856
rect 77502 2 78530 856
rect 78698 2 79634 856
rect 79802 2 80830 856
rect 80998 2 82026 856
rect 82194 2 83222 856
rect 83390 2 84418 856
rect 84586 2 85614 856
rect 85782 2 86810 856
rect 86978 2 87914 856
rect 88082 2 89110 856
rect 89278 2 90306 856
rect 90474 2 91502 856
rect 91670 2 92698 856
rect 92866 2 93894 856
rect 94062 2 95090 856
rect 95258 2 96194 856
rect 96362 2 97390 856
rect 97558 2 98586 856
rect 98754 2 99782 856
rect 99950 2 100978 856
rect 101146 2 102174 856
rect 102342 2 103278 856
rect 103446 2 104474 856
rect 104642 2 105670 856
rect 105838 2 106866 856
rect 107034 2 108062 856
rect 108230 2 109258 856
rect 109426 2 110454 856
rect 110622 2 111558 856
rect 111726 2 112754 856
rect 112922 2 113950 856
rect 114118 2 115146 856
rect 115314 2 116342 856
rect 116510 2 117538 856
rect 117706 2 118734 856
rect 118902 2 119838 856
rect 120006 2 121034 856
rect 121202 2 122230 856
rect 122398 2 123426 856
rect 123594 2 124622 856
rect 124790 2 125818 856
rect 125986 2 126922 856
rect 127090 2 128118 856
rect 128286 2 129314 856
rect 129482 2 130510 856
rect 130678 2 131706 856
rect 131874 2 132902 856
rect 133070 2 134098 856
rect 134266 2 135202 856
rect 135370 2 136398 856
rect 136566 2 137594 856
rect 137762 2 138790 856
rect 138958 2 139986 856
rect 140154 2 141182 856
rect 141350 2 142378 856
rect 142546 2 143482 856
rect 143650 2 144678 856
rect 144846 2 145874 856
rect 146042 2 147070 856
rect 147238 2 148266 856
rect 148434 2 149462 856
rect 149630 2 150566 856
rect 150734 2 151762 856
rect 151930 2 152958 856
rect 153126 2 154154 856
rect 154322 2 155350 856
rect 155518 2 156546 856
rect 156714 2 157742 856
rect 157910 2 158846 856
rect 159014 2 160042 856
rect 160210 2 161238 856
rect 161406 2 162434 856
rect 162602 2 163630 856
rect 163798 2 164826 856
rect 164994 2 166022 856
rect 166190 2 167126 856
rect 167294 2 168322 856
rect 168490 2 169518 856
rect 169686 2 170714 856
rect 170882 2 171910 856
rect 172078 2 173106 856
rect 173274 2 174210 856
rect 174378 2 175406 856
rect 175574 2 176602 856
rect 176770 2 177798 856
rect 177966 2 178994 856
rect 179162 2 180190 856
rect 180358 2 181386 856
rect 181554 2 182490 856
rect 182658 2 183686 856
rect 183854 2 184882 856
rect 185050 2 186078 856
rect 186246 2 187274 856
rect 187442 2 188470 856
rect 188638 2 189666 856
rect 189834 2 190770 856
rect 190938 2 191966 856
rect 192134 2 193162 856
rect 193330 2 194358 856
rect 194526 2 195554 856
rect 195722 2 196750 856
rect 196918 2 197854 856
rect 198022 2 199050 856
rect 199218 2 200246 856
rect 200414 2 201442 856
rect 201610 2 202638 856
rect 202806 2 203834 856
rect 204002 2 205030 856
rect 205198 2 206134 856
rect 206302 2 207330 856
rect 207498 2 208526 856
rect 208694 2 209722 856
rect 209890 2 210918 856
rect 211086 2 212114 856
rect 212282 2 213310 856
rect 213478 2 214414 856
rect 214582 2 215610 856
rect 215778 2 216806 856
rect 216974 2 218002 856
rect 218170 2 219198 856
rect 219366 2 220394 856
rect 220562 2 221498 856
rect 221666 2 222694 856
rect 222862 2 223890 856
rect 224058 2 225086 856
rect 225254 2 226282 856
rect 226450 2 227478 856
rect 227646 2 228674 856
rect 228842 2 229778 856
rect 229946 2 230974 856
rect 231142 2 232170 856
rect 232338 2 233366 856
rect 233534 2 234562 856
rect 234730 2 235758 856
rect 235926 2 236954 856
rect 237122 2 238058 856
rect 238226 2 239254 856
rect 239422 2 240450 856
rect 240618 2 241646 856
rect 241814 2 242842 856
rect 243010 2 244038 856
rect 244206 2 245142 856
rect 245310 2 246338 856
rect 246506 2 247534 856
rect 247702 2 248730 856
rect 248898 2 249926 856
rect 250094 2 251122 856
rect 251290 2 252318 856
rect 252486 2 253422 856
rect 253590 2 254618 856
rect 254786 2 255814 856
rect 255982 2 257010 856
rect 257178 2 258206 856
rect 258374 2 259402 856
rect 259570 2 260598 856
rect 260766 2 261702 856
rect 261870 2 262898 856
rect 263066 2 264094 856
rect 264262 2 265290 856
rect 265458 2 266486 856
rect 266654 2 267682 856
rect 267850 2 268786 856
rect 268954 2 269982 856
rect 270150 2 271178 856
rect 271346 2 272374 856
rect 272542 2 273570 856
rect 273738 2 274766 856
rect 274934 2 275962 856
rect 276130 2 277066 856
rect 277234 2 278262 856
rect 278430 2 279458 856
rect 279626 2 280654 856
rect 280822 2 281850 856
rect 282018 2 283046 856
rect 283214 2 284242 856
rect 284410 2 285346 856
rect 285514 2 286542 856
rect 286710 2 287738 856
rect 287906 2 288934 856
rect 289102 2 290130 856
rect 290298 2 291326 856
rect 291494 2 292522 856
rect 292690 2 293626 856
rect 293794 2 294822 856
rect 294990 2 296018 856
rect 296186 2 297214 856
rect 297382 2 298410 856
rect 298578 2 299606 856
rect 299774 2 300710 856
rect 300878 2 301906 856
rect 302074 2 303102 856
rect 303270 2 304298 856
rect 304466 2 305494 856
rect 305662 2 306690 856
rect 306858 2 307886 856
rect 308054 2 308990 856
rect 309158 2 310186 856
rect 310354 2 311382 856
rect 311550 2 312578 856
rect 312746 2 313774 856
rect 313942 2 314970 856
rect 315138 2 316166 856
rect 316334 2 317270 856
rect 317438 2 318466 856
rect 318634 2 319662 856
rect 319830 2 320858 856
rect 321026 2 322054 856
rect 322222 2 323250 856
rect 323418 2 324354 856
rect 324522 2 325550 856
rect 325718 2 326746 856
rect 326914 2 327942 856
rect 328110 2 329138 856
rect 329306 2 330334 856
rect 330502 2 331530 856
rect 331698 2 332634 856
rect 332802 2 333830 856
rect 333998 2 335026 856
rect 335194 2 336222 856
rect 336390 2 337418 856
rect 337586 2 338614 856
rect 338782 2 339810 856
rect 339978 2 340914 856
rect 341082 2 342110 856
rect 342278 2 343306 856
rect 343474 2 344502 856
rect 344670 2 345698 856
rect 345866 2 346894 856
rect 347062 2 347998 856
rect 348166 2 349194 856
rect 349362 2 350390 856
rect 350558 2 351586 856
rect 351754 2 352782 856
rect 352950 2 353978 856
rect 354146 2 355174 856
rect 355342 2 356278 856
rect 356446 2 357474 856
rect 357642 2 358670 856
rect 358838 2 359866 856
rect 360034 2 361062 856
rect 361230 2 362258 856
rect 362426 2 363454 856
rect 363622 2 364558 856
rect 364726 2 365754 856
rect 365922 2 366950 856
rect 367118 2 368146 856
rect 368314 2 369342 856
rect 369510 2 370538 856
rect 370706 2 371642 856
rect 371810 2 372838 856
rect 373006 2 374034 856
rect 374202 2 375230 856
rect 375398 2 376426 856
rect 376594 2 377622 856
rect 377790 2 378818 856
rect 378986 2 379922 856
rect 380090 2 381118 856
rect 381286 2 382314 856
rect 382482 2 383510 856
rect 383678 2 384706 856
rect 384874 2 385902 856
rect 386070 2 387098 856
rect 387266 2 388202 856
rect 388370 2 389398 856
rect 389566 2 390594 856
rect 390762 2 391790 856
rect 391958 2 392986 856
rect 393154 2 394182 856
rect 394350 2 395286 856
rect 395454 2 396482 856
rect 396650 2 397678 856
rect 397846 2 398874 856
rect 399042 2 400070 856
rect 400238 2 401266 856
rect 401434 2 402462 856
rect 402630 2 403566 856
rect 403734 2 404762 856
rect 404930 2 405958 856
rect 406126 2 407154 856
rect 407322 2 408350 856
rect 408518 2 409546 856
rect 409714 2 410742 856
rect 410910 2 411846 856
rect 412014 2 413042 856
rect 413210 2 414238 856
rect 414406 2 415434 856
rect 415602 2 416630 856
rect 416798 2 417826 856
rect 417994 2 418930 856
rect 419098 2 420126 856
rect 420294 2 421322 856
rect 421490 2 422518 856
rect 422686 2 423714 856
rect 423882 2 424910 856
rect 425078 2 426106 856
rect 426274 2 427210 856
rect 427378 2 428406 856
rect 428574 2 429602 856
rect 429770 2 430798 856
rect 430966 2 431994 856
rect 432162 2 433190 856
rect 433358 2 434386 856
rect 434554 2 435490 856
rect 435658 2 436686 856
rect 436854 2 437882 856
rect 438050 2 439078 856
rect 439246 2 440274 856
rect 440442 2 441470 856
rect 441638 2 442574 856
rect 442742 2 443770 856
rect 443938 2 444966 856
rect 445134 2 446162 856
rect 446330 2 447358 856
rect 447526 2 448554 856
rect 448722 2 449750 856
rect 449918 2 450854 856
rect 451022 2 452050 856
rect 452218 2 453246 856
rect 453414 2 454442 856
rect 454610 2 455638 856
rect 455806 2 456834 856
rect 457002 2 458030 856
rect 458198 2 459134 856
rect 459302 2 460330 856
rect 460498 2 461526 856
rect 461694 2 462722 856
rect 462890 2 463918 856
rect 464086 2 465114 856
rect 465282 2 466218 856
rect 466386 2 467414 856
rect 467582 2 468610 856
rect 468778 2 469806 856
rect 469974 2 471002 856
rect 471170 2 472198 856
rect 472366 2 473394 856
rect 473562 2 474498 856
rect 474666 2 475694 856
rect 475862 2 476890 856
rect 477058 2 478086 856
rect 478254 2 479282 856
rect 479450 2 480478 856
rect 480646 2 481674 856
rect 481842 2 482778 856
rect 482946 2 483974 856
rect 484142 2 485170 856
rect 485338 2 486366 856
rect 486534 2 487562 856
rect 487730 2 488758 856
rect 488926 2 489862 856
rect 490030 2 491058 856
rect 491226 2 492254 856
rect 492422 2 493450 856
rect 493618 2 494646 856
rect 494814 2 495842 856
rect 496010 2 497038 856
rect 497206 2 498142 856
rect 498310 2 499338 856
rect 499506 2 500534 856
rect 500702 2 501730 856
rect 501898 2 502926 856
rect 503094 2 504122 856
rect 504290 2 505318 856
rect 505486 2 506422 856
rect 506590 2 507618 856
rect 507786 2 508814 856
rect 508982 2 510010 856
rect 510178 2 511206 856
rect 511374 2 512402 856
rect 512570 2 513506 856
rect 513674 2 514702 856
rect 514870 2 515898 856
rect 516066 2 517094 856
rect 517262 2 518290 856
rect 518458 2 519486 856
rect 519654 2 520682 856
rect 520850 2 521786 856
rect 521954 2 522982 856
rect 523150 2 524178 856
rect 524346 2 525374 856
rect 525542 2 526570 856
rect 526738 2 527766 856
rect 527934 2 528962 856
rect 529130 2 530066 856
rect 530234 2 531262 856
rect 531430 2 532458 856
rect 532626 2 533654 856
rect 533822 2 534850 856
rect 535018 2 536046 856
rect 536214 2 537150 856
rect 537318 2 538346 856
rect 538514 2 539542 856
rect 539710 2 540738 856
rect 540906 2 541934 856
rect 542102 2 543130 856
rect 543298 2 544326 856
rect 544494 2 545430 856
rect 545598 2 546626 856
rect 546794 2 547822 856
rect 547990 2 549018 856
rect 549186 2 550214 856
rect 550382 2 551410 856
rect 551578 2 552606 856
rect 552774 2 553710 856
rect 553878 2 554906 856
rect 555074 2 556102 856
rect 556270 2 557298 856
rect 557466 2 558494 856
rect 558662 2 559690 856
rect 559858 2 560794 856
rect 560962 2 561990 856
rect 562158 2 563186 856
rect 563354 2 564382 856
rect 564550 2 565578 856
rect 565746 2 566774 856
rect 566942 2 567970 856
rect 568138 2 569074 856
rect 569242 2 570270 856
rect 570438 2 571466 856
rect 571634 2 572662 856
rect 572830 2 573858 856
rect 574026 2 575054 856
rect 575222 2 576250 856
rect 576418 2 577354 856
rect 577522 2 578550 856
rect 578718 2 579746 856
rect 579914 2 580942 856
rect 581110 2 582138 856
rect 582306 2 583334 856
<< metal3 >>
rect 0 697280 800 697400
rect 583200 697144 584000 697264
rect 0 684224 800 684344
rect 583200 683816 584000 683936
rect 0 671168 800 671288
rect 583200 670624 584000 670744
rect 0 658112 800 658232
rect 583200 657296 584000 657416
rect 0 645056 800 645176
rect 583200 643968 584000 644088
rect 0 632000 800 632120
rect 583200 630776 584000 630896
rect 0 619080 800 619200
rect 583200 617448 584000 617568
rect 0 606024 800 606144
rect 583200 604120 584000 604240
rect 0 592968 800 593088
rect 583200 590928 584000 591048
rect 0 579912 800 580032
rect 583200 577600 584000 577720
rect 0 566856 800 566976
rect 583200 564272 584000 564392
rect 0 553800 800 553920
rect 583200 551080 584000 551200
rect 0 540744 800 540864
rect 583200 537752 584000 537872
rect 0 527824 800 527944
rect 583200 524424 584000 524544
rect 0 514768 800 514888
rect 583200 511232 584000 511352
rect 0 501712 800 501832
rect 583200 497904 584000 498024
rect 0 488656 800 488776
rect 583200 484576 584000 484696
rect 0 475600 800 475720
rect 583200 471384 584000 471504
rect 0 462544 800 462664
rect 583200 458056 584000 458176
rect 0 449488 800 449608
rect 583200 444728 584000 444848
rect 0 436568 800 436688
rect 583200 431536 584000 431656
rect 0 423512 800 423632
rect 583200 418208 584000 418328
rect 0 410456 800 410576
rect 583200 404880 584000 405000
rect 0 397400 800 397520
rect 583200 391688 584000 391808
rect 0 384344 800 384464
rect 583200 378360 584000 378480
rect 0 371288 800 371408
rect 583200 365032 584000 365152
rect 0 358368 800 358488
rect 583200 351840 584000 351960
rect 0 345312 800 345432
rect 583200 338512 584000 338632
rect 0 332256 800 332376
rect 583200 325184 584000 325304
rect 0 319200 800 319320
rect 583200 311992 584000 312112
rect 0 306144 800 306264
rect 583200 298664 584000 298784
rect 0 293088 800 293208
rect 583200 285336 584000 285456
rect 0 280032 800 280152
rect 583200 272144 584000 272264
rect 0 267112 800 267232
rect 583200 258816 584000 258936
rect 0 254056 800 254176
rect 583200 245488 584000 245608
rect 0 241000 800 241120
rect 583200 232296 584000 232416
rect 0 227944 800 228064
rect 583200 218968 584000 219088
rect 0 214888 800 215008
rect 583200 205640 584000 205760
rect 0 201832 800 201952
rect 583200 192448 584000 192568
rect 0 188776 800 188896
rect 583200 179120 584000 179240
rect 0 175856 800 175976
rect 583200 165792 584000 165912
rect 0 162800 800 162920
rect 583200 152600 584000 152720
rect 0 149744 800 149864
rect 583200 139272 584000 139392
rect 0 136688 800 136808
rect 583200 125944 584000 126064
rect 0 123632 800 123752
rect 583200 112752 584000 112872
rect 0 110576 800 110696
rect 583200 99424 584000 99544
rect 0 97520 800 97640
rect 583200 86096 584000 86216
rect 0 84600 800 84720
rect 583200 72904 584000 73024
rect 0 71544 800 71664
rect 583200 59576 584000 59696
rect 0 58488 800 58608
rect 583200 46248 584000 46368
rect 0 45432 800 45552
rect 583200 33056 584000 33176
rect 0 32376 800 32496
rect 583200 19728 584000 19848
rect 0 19320 800 19440
rect 0 6400 800 6520
rect 583200 6536 584000 6656
<< obsm3 >>
rect 800 697480 583200 701793
rect 880 697344 583200 697480
rect 880 697200 583120 697344
rect 800 697064 583120 697200
rect 800 684424 583200 697064
rect 880 684144 583200 684424
rect 800 684016 583200 684144
rect 800 683736 583120 684016
rect 800 671368 583200 683736
rect 880 671088 583200 671368
rect 800 670824 583200 671088
rect 800 670544 583120 670824
rect 800 658312 583200 670544
rect 880 658032 583200 658312
rect 800 657496 583200 658032
rect 800 657216 583120 657496
rect 800 645256 583200 657216
rect 880 644976 583200 645256
rect 800 644168 583200 644976
rect 800 643888 583120 644168
rect 800 632200 583200 643888
rect 880 631920 583200 632200
rect 800 630976 583200 631920
rect 800 630696 583120 630976
rect 800 619280 583200 630696
rect 880 619000 583200 619280
rect 800 617648 583200 619000
rect 800 617368 583120 617648
rect 800 606224 583200 617368
rect 880 605944 583200 606224
rect 800 604320 583200 605944
rect 800 604040 583120 604320
rect 800 593168 583200 604040
rect 880 592888 583200 593168
rect 800 591128 583200 592888
rect 800 590848 583120 591128
rect 800 580112 583200 590848
rect 880 579832 583200 580112
rect 800 577800 583200 579832
rect 800 577520 583120 577800
rect 800 567056 583200 577520
rect 880 566776 583200 567056
rect 800 564472 583200 566776
rect 800 564192 583120 564472
rect 800 554000 583200 564192
rect 880 553720 583200 554000
rect 800 551280 583200 553720
rect 800 551000 583120 551280
rect 800 540944 583200 551000
rect 880 540664 583200 540944
rect 800 537952 583200 540664
rect 800 537672 583120 537952
rect 800 528024 583200 537672
rect 880 527744 583200 528024
rect 800 524624 583200 527744
rect 800 524344 583120 524624
rect 800 514968 583200 524344
rect 880 514688 583200 514968
rect 800 511432 583200 514688
rect 800 511152 583120 511432
rect 800 501912 583200 511152
rect 880 501632 583200 501912
rect 800 498104 583200 501632
rect 800 497824 583120 498104
rect 800 488856 583200 497824
rect 880 488576 583200 488856
rect 800 484776 583200 488576
rect 800 484496 583120 484776
rect 800 475800 583200 484496
rect 880 475520 583200 475800
rect 800 471584 583200 475520
rect 800 471304 583120 471584
rect 800 462744 583200 471304
rect 880 462464 583200 462744
rect 800 458256 583200 462464
rect 800 457976 583120 458256
rect 800 449688 583200 457976
rect 880 449408 583200 449688
rect 800 444928 583200 449408
rect 800 444648 583120 444928
rect 800 436768 583200 444648
rect 880 436488 583200 436768
rect 800 431736 583200 436488
rect 800 431456 583120 431736
rect 800 423712 583200 431456
rect 880 423432 583200 423712
rect 800 418408 583200 423432
rect 800 418128 583120 418408
rect 800 410656 583200 418128
rect 880 410376 583200 410656
rect 800 405080 583200 410376
rect 800 404800 583120 405080
rect 800 397600 583200 404800
rect 880 397320 583200 397600
rect 800 391888 583200 397320
rect 800 391608 583120 391888
rect 800 384544 583200 391608
rect 880 384264 583200 384544
rect 800 378560 583200 384264
rect 800 378280 583120 378560
rect 800 371488 583200 378280
rect 880 371208 583200 371488
rect 800 365232 583200 371208
rect 800 364952 583120 365232
rect 800 358568 583200 364952
rect 880 358288 583200 358568
rect 800 352040 583200 358288
rect 800 351760 583120 352040
rect 800 345512 583200 351760
rect 880 345232 583200 345512
rect 800 338712 583200 345232
rect 800 338432 583120 338712
rect 800 332456 583200 338432
rect 880 332176 583200 332456
rect 800 325384 583200 332176
rect 800 325104 583120 325384
rect 800 319400 583200 325104
rect 880 319120 583200 319400
rect 800 312192 583200 319120
rect 800 311912 583120 312192
rect 800 306344 583200 311912
rect 880 306064 583200 306344
rect 800 298864 583200 306064
rect 800 298584 583120 298864
rect 800 293288 583200 298584
rect 880 293008 583200 293288
rect 800 285536 583200 293008
rect 800 285256 583120 285536
rect 800 280232 583200 285256
rect 880 279952 583200 280232
rect 800 272344 583200 279952
rect 800 272064 583120 272344
rect 800 267312 583200 272064
rect 880 267032 583200 267312
rect 800 259016 583200 267032
rect 800 258736 583120 259016
rect 800 254256 583200 258736
rect 880 253976 583200 254256
rect 800 245688 583200 253976
rect 800 245408 583120 245688
rect 800 241200 583200 245408
rect 880 240920 583200 241200
rect 800 232496 583200 240920
rect 800 232216 583120 232496
rect 800 228144 583200 232216
rect 880 227864 583200 228144
rect 800 219168 583200 227864
rect 800 218888 583120 219168
rect 800 215088 583200 218888
rect 880 214808 583200 215088
rect 800 205840 583200 214808
rect 800 205560 583120 205840
rect 800 202032 583200 205560
rect 880 201752 583200 202032
rect 800 192648 583200 201752
rect 800 192368 583120 192648
rect 800 188976 583200 192368
rect 880 188696 583200 188976
rect 800 179320 583200 188696
rect 800 179040 583120 179320
rect 800 176056 583200 179040
rect 880 175776 583200 176056
rect 800 165992 583200 175776
rect 800 165712 583120 165992
rect 800 163000 583200 165712
rect 880 162720 583200 163000
rect 800 152800 583200 162720
rect 800 152520 583120 152800
rect 800 149944 583200 152520
rect 880 149664 583200 149944
rect 800 139472 583200 149664
rect 800 139192 583120 139472
rect 800 136888 583200 139192
rect 880 136608 583200 136888
rect 800 126144 583200 136608
rect 800 125864 583120 126144
rect 800 123832 583200 125864
rect 880 123552 583200 123832
rect 800 112952 583200 123552
rect 800 112672 583120 112952
rect 800 110776 583200 112672
rect 880 110496 583200 110776
rect 800 99624 583200 110496
rect 800 99344 583120 99624
rect 800 97720 583200 99344
rect 880 97440 583200 97720
rect 800 86296 583200 97440
rect 800 86016 583120 86296
rect 800 84800 583200 86016
rect 880 84520 583200 84800
rect 800 73104 583200 84520
rect 800 72824 583120 73104
rect 800 71744 583200 72824
rect 880 71464 583200 71744
rect 800 59776 583200 71464
rect 800 59496 583120 59776
rect 800 58688 583200 59496
rect 880 58408 583200 58688
rect 800 46448 583200 58408
rect 800 46168 583120 46448
rect 800 45632 583200 46168
rect 880 45352 583200 45632
rect 800 33256 583200 45352
rect 800 32976 583120 33256
rect 800 32576 583200 32976
rect 880 32296 583200 32576
rect 800 19928 583200 32296
rect 800 19648 583120 19928
rect 800 19520 583200 19648
rect 880 19240 583200 19520
rect 800 6736 583200 19240
rect 800 6600 583120 6736
rect 880 6456 583120 6600
rect 880 6320 583200 6456
rect 800 1259 583200 6320
<< metal4 >>
rect -916 156 -596 703780
rect -256 816 64 703120
rect 5944 156 6264 703780
rect 12944 156 13264 703780
rect 19944 653408 20264 703780
rect 26944 653408 27264 703780
rect 33944 653408 34264 703780
rect 40944 653408 41264 703780
rect 47944 653408 48264 703780
rect 54944 653408 55264 703780
rect 19944 597408 20264 608048
rect 26944 597408 27264 608048
rect 33944 597408 34264 608048
rect 40944 597408 41264 608048
rect 47944 597408 48264 608048
rect 54944 597408 55264 608048
rect 19944 541408 20264 552048
rect 26944 541408 27264 552048
rect 33944 541408 34264 552048
rect 40944 541408 41264 552048
rect 47944 541408 48264 552048
rect 54944 541408 55264 552048
rect 19944 485408 20264 496048
rect 26944 485408 27264 496048
rect 33944 485408 34264 496048
rect 40944 485408 41264 496048
rect 47944 485408 48264 496048
rect 54944 485408 55264 496048
rect 19944 429408 20264 440048
rect 26944 429408 27264 440048
rect 33944 429408 34264 440048
rect 40944 429408 41264 440048
rect 47944 429408 48264 440048
rect 54944 429408 55264 440048
rect 19944 373408 20264 384048
rect 26944 373408 27264 384048
rect 33944 373408 34264 384048
rect 40944 373408 41264 384048
rect 47944 373408 48264 384048
rect 54944 373408 55264 384048
rect 19944 317408 20264 328048
rect 26944 317408 27264 328048
rect 33944 317408 34264 328048
rect 40944 317408 41264 328048
rect 47944 317408 48264 328048
rect 54944 317408 55264 328048
rect 19944 261408 20264 272048
rect 26944 261408 27264 272048
rect 33944 261408 34264 272048
rect 40944 261408 41264 272048
rect 47944 261408 48264 272048
rect 54944 261408 55264 272048
rect 19944 205408 20264 216048
rect 26944 205408 27264 216048
rect 33944 205408 34264 216048
rect 40944 205408 41264 216048
rect 47944 205408 48264 216048
rect 54944 205408 55264 216048
rect 19944 149408 20264 160048
rect 26944 149408 27264 160048
rect 33944 149408 34264 160048
rect 40944 149408 41264 160048
rect 47944 149408 48264 160048
rect 54944 149408 55264 160048
rect 19944 93408 20264 104048
rect 26944 93408 27264 104048
rect 33944 93408 34264 104048
rect 40944 93408 41264 104048
rect 47944 93408 48264 104048
rect 54944 93408 55264 104048
rect 19944 156 20264 48048
rect 26944 156 27264 48048
rect 33944 156 34264 48048
rect 40944 156 41264 48048
rect 47944 156 48264 48048
rect 54944 156 55264 48048
rect 61944 156 62264 703780
rect 68944 156 69264 703780
rect 75944 653408 76264 703780
rect 82944 653408 83264 703780
rect 89944 653408 90264 703780
rect 96944 653408 97264 703780
rect 103944 653408 104264 703780
rect 110944 653408 111264 703780
rect 75944 597408 76264 608048
rect 82944 597408 83264 608048
rect 89944 597408 90264 608048
rect 96944 597408 97264 608048
rect 103944 597408 104264 608048
rect 110944 597408 111264 608048
rect 75944 541408 76264 552048
rect 82944 541408 83264 552048
rect 89944 541408 90264 552048
rect 96944 541408 97264 552048
rect 103944 541408 104264 552048
rect 110944 541408 111264 552048
rect 75944 485408 76264 496048
rect 82944 485408 83264 496048
rect 89944 485408 90264 496048
rect 96944 485408 97264 496048
rect 103944 485408 104264 496048
rect 110944 485408 111264 496048
rect 75944 429408 76264 440048
rect 82944 429408 83264 440048
rect 89944 429408 90264 440048
rect 96944 429408 97264 440048
rect 103944 429408 104264 440048
rect 110944 429408 111264 440048
rect 75944 373408 76264 384048
rect 82944 373408 83264 384048
rect 89944 373408 90264 384048
rect 96944 373408 97264 384048
rect 103944 373408 104264 384048
rect 110944 373408 111264 384048
rect 75944 317408 76264 328048
rect 82944 317408 83264 328048
rect 89944 317408 90264 328048
rect 96944 317408 97264 328048
rect 103944 317408 104264 328048
rect 110944 317408 111264 328048
rect 75944 261408 76264 272048
rect 82944 261408 83264 272048
rect 89944 261408 90264 272048
rect 96944 261408 97264 272048
rect 103944 261408 104264 272048
rect 110944 261408 111264 272048
rect 75944 205408 76264 216048
rect 82944 205408 83264 216048
rect 89944 205408 90264 216048
rect 96944 205408 97264 216048
rect 103944 205408 104264 216048
rect 110944 205408 111264 216048
rect 75944 149408 76264 160048
rect 82944 149408 83264 160048
rect 89944 149408 90264 160048
rect 96944 149408 97264 160048
rect 103944 149408 104264 160048
rect 110944 149408 111264 160048
rect 75944 93408 76264 104048
rect 82944 93408 83264 104048
rect 89944 93408 90264 104048
rect 96944 93408 97264 104048
rect 103944 93408 104264 104048
rect 110944 93408 111264 104048
rect 75944 156 76264 48048
rect 82944 156 83264 48048
rect 89944 156 90264 48048
rect 96944 156 97264 48048
rect 103944 156 104264 48048
rect 110944 156 111264 48048
rect 117944 156 118264 703780
rect 124944 156 125264 703780
rect 131944 653408 132264 703780
rect 138944 653408 139264 703780
rect 145944 653408 146264 703780
rect 152944 653408 153264 703780
rect 159944 653408 160264 703780
rect 166944 653408 167264 703780
rect 131944 597408 132264 608048
rect 138944 597408 139264 608048
rect 145944 597408 146264 608048
rect 152944 597408 153264 608048
rect 159944 597408 160264 608048
rect 166944 597408 167264 608048
rect 131944 541408 132264 552048
rect 138944 541408 139264 552048
rect 145944 541408 146264 552048
rect 152944 541408 153264 552048
rect 159944 541408 160264 552048
rect 166944 541408 167264 552048
rect 131944 485408 132264 496048
rect 138944 485408 139264 496048
rect 145944 485408 146264 496048
rect 152944 485408 153264 496048
rect 159944 485408 160264 496048
rect 166944 485408 167264 496048
rect 131944 429408 132264 440048
rect 138944 429408 139264 440048
rect 145944 429408 146264 440048
rect 152944 429408 153264 440048
rect 159944 429408 160264 440048
rect 166944 429408 167264 440048
rect 131944 373408 132264 384048
rect 138944 373408 139264 384048
rect 145944 373408 146264 384048
rect 152944 373408 153264 384048
rect 159944 373408 160264 384048
rect 166944 373408 167264 384048
rect 131944 317408 132264 328048
rect 138944 317408 139264 328048
rect 145944 317408 146264 328048
rect 152944 317408 153264 328048
rect 159944 317408 160264 328048
rect 166944 317408 167264 328048
rect 131944 261408 132264 272048
rect 138944 261408 139264 272048
rect 145944 261408 146264 272048
rect 152944 261408 153264 272048
rect 159944 261408 160264 272048
rect 166944 261408 167264 272048
rect 131944 205408 132264 216048
rect 138944 205408 139264 216048
rect 145944 205408 146264 216048
rect 152944 205408 153264 216048
rect 159944 205408 160264 216048
rect 166944 205408 167264 216048
rect 131944 149408 132264 160048
rect 138944 149408 139264 160048
rect 145944 149408 146264 160048
rect 152944 149408 153264 160048
rect 159944 149408 160264 160048
rect 166944 149408 167264 160048
rect 131944 93408 132264 104048
rect 138944 93408 139264 104048
rect 145944 93408 146264 104048
rect 152944 93408 153264 104048
rect 159944 93408 160264 104048
rect 166944 93408 167264 104048
rect 131944 156 132264 48048
rect 138944 156 139264 48048
rect 145944 156 146264 48048
rect 152944 156 153264 48048
rect 159944 156 160264 48048
rect 166944 156 167264 48048
rect 173944 156 174264 703780
rect 180944 156 181264 703780
rect 187944 653408 188264 703780
rect 194944 653408 195264 703780
rect 201944 653408 202264 703780
rect 208944 653408 209264 703780
rect 215944 653408 216264 703780
rect 222944 653408 223264 703780
rect 187944 597408 188264 608048
rect 194944 597408 195264 608048
rect 201944 597408 202264 608048
rect 208944 597408 209264 608048
rect 215944 597408 216264 608048
rect 222944 597408 223264 608048
rect 187944 541408 188264 552048
rect 194944 541408 195264 552048
rect 201944 541408 202264 552048
rect 208944 541408 209264 552048
rect 215944 541408 216264 552048
rect 222944 541408 223264 552048
rect 187944 485408 188264 496048
rect 194944 485408 195264 496048
rect 201944 485408 202264 496048
rect 208944 485408 209264 496048
rect 215944 485408 216264 496048
rect 222944 485408 223264 496048
rect 187944 429408 188264 440048
rect 194944 429408 195264 440048
rect 201944 429408 202264 440048
rect 208944 429408 209264 440048
rect 215944 429408 216264 440048
rect 222944 429408 223264 440048
rect 187944 373408 188264 384048
rect 194944 373408 195264 384048
rect 201944 373408 202264 384048
rect 208944 373408 209264 384048
rect 215944 373408 216264 384048
rect 222944 373408 223264 384048
rect 187944 317408 188264 328048
rect 194944 317408 195264 328048
rect 201944 317408 202264 328048
rect 208944 317408 209264 328048
rect 215944 317408 216264 328048
rect 222944 317408 223264 328048
rect 187944 261408 188264 272048
rect 194944 261408 195264 272048
rect 201944 261408 202264 272048
rect 208944 261408 209264 272048
rect 215944 261408 216264 272048
rect 222944 261408 223264 272048
rect 187944 205408 188264 216048
rect 194944 205408 195264 216048
rect 201944 205408 202264 216048
rect 208944 205408 209264 216048
rect 215944 205408 216264 216048
rect 222944 205408 223264 216048
rect 187944 149408 188264 160048
rect 194944 149408 195264 160048
rect 201944 149408 202264 160048
rect 208944 149408 209264 160048
rect 215944 149408 216264 160048
rect 222944 149408 223264 160048
rect 187944 93408 188264 104048
rect 194944 93408 195264 104048
rect 201944 93408 202264 104048
rect 208944 93408 209264 104048
rect 215944 93408 216264 104048
rect 222944 93408 223264 104048
rect 187944 156 188264 48048
rect 194944 156 195264 48048
rect 201944 156 202264 48048
rect 208944 156 209264 48048
rect 215944 156 216264 48048
rect 222944 156 223264 48048
rect 229944 156 230264 703780
rect 236944 156 237264 703780
rect 243944 653408 244264 703780
rect 250944 653408 251264 703780
rect 257944 653408 258264 703780
rect 264944 653408 265264 703780
rect 271944 653408 272264 703780
rect 278944 653408 279264 703780
rect 243944 597408 244264 608048
rect 250944 597408 251264 608048
rect 257944 597408 258264 608048
rect 264944 597408 265264 608048
rect 271944 597408 272264 608048
rect 278944 597408 279264 608048
rect 243944 541408 244264 552048
rect 250944 541408 251264 552048
rect 257944 541408 258264 552048
rect 264944 541408 265264 552048
rect 271944 541408 272264 552048
rect 278944 541408 279264 552048
rect 243944 485408 244264 496048
rect 250944 485408 251264 496048
rect 257944 485408 258264 496048
rect 264944 485408 265264 496048
rect 271944 485408 272264 496048
rect 278944 485408 279264 496048
rect 243944 429408 244264 440048
rect 250944 429408 251264 440048
rect 257944 429408 258264 440048
rect 264944 429408 265264 440048
rect 271944 429408 272264 440048
rect 278944 429408 279264 440048
rect 243944 373408 244264 384048
rect 250944 373408 251264 384048
rect 257944 373408 258264 384048
rect 264944 373408 265264 384048
rect 271944 373408 272264 384048
rect 278944 373408 279264 384048
rect 243944 317408 244264 328048
rect 250944 317408 251264 328048
rect 257944 317408 258264 328048
rect 264944 317408 265264 328048
rect 271944 317408 272264 328048
rect 278944 317408 279264 328048
rect 243944 261408 244264 272048
rect 250944 261408 251264 272048
rect 257944 261408 258264 272048
rect 264944 261408 265264 272048
rect 271944 261408 272264 272048
rect 278944 261408 279264 272048
rect 243944 205408 244264 216048
rect 250944 205408 251264 216048
rect 257944 205408 258264 216048
rect 264944 205408 265264 216048
rect 271944 205408 272264 216048
rect 278944 205408 279264 216048
rect 243944 149408 244264 160048
rect 250944 149408 251264 160048
rect 257944 149408 258264 160048
rect 264944 149408 265264 160048
rect 271944 149408 272264 160048
rect 278944 149408 279264 160048
rect 243944 93408 244264 104048
rect 250944 93408 251264 104048
rect 257944 93408 258264 104048
rect 264944 93408 265264 104048
rect 271944 93408 272264 104048
rect 278944 93408 279264 104048
rect 243944 156 244264 48048
rect 250944 156 251264 48048
rect 257944 156 258264 48048
rect 264944 156 265264 48048
rect 271944 156 272264 48048
rect 278944 156 279264 48048
rect 285944 156 286264 703780
rect 292944 156 293264 703780
rect 299944 653408 300264 703780
rect 306944 653408 307264 703780
rect 313944 653408 314264 703780
rect 320944 653408 321264 703780
rect 327944 653408 328264 703780
rect 334944 653408 335264 703780
rect 299944 597408 300264 608048
rect 306944 597408 307264 608048
rect 313944 597408 314264 608048
rect 320944 597408 321264 608048
rect 327944 597408 328264 608048
rect 334944 597408 335264 608048
rect 299944 541408 300264 552048
rect 306944 541408 307264 552048
rect 313944 541408 314264 552048
rect 320944 541408 321264 552048
rect 327944 541408 328264 552048
rect 334944 541408 335264 552048
rect 299944 485408 300264 496048
rect 306944 485408 307264 496048
rect 313944 485408 314264 496048
rect 320944 485408 321264 496048
rect 327944 485408 328264 496048
rect 334944 485408 335264 496048
rect 299944 429408 300264 440048
rect 306944 429408 307264 440048
rect 313944 429408 314264 440048
rect 320944 429408 321264 440048
rect 327944 429408 328264 440048
rect 334944 429408 335264 440048
rect 299944 373408 300264 384048
rect 306944 373408 307264 384048
rect 313944 373408 314264 384048
rect 320944 373408 321264 384048
rect 327944 373408 328264 384048
rect 334944 373408 335264 384048
rect 299944 317408 300264 328048
rect 306944 317408 307264 328048
rect 313944 317408 314264 328048
rect 320944 317408 321264 328048
rect 327944 317408 328264 328048
rect 334944 317408 335264 328048
rect 299944 261408 300264 272048
rect 306944 261408 307264 272048
rect 313944 261408 314264 272048
rect 320944 261408 321264 272048
rect 327944 261408 328264 272048
rect 334944 261408 335264 272048
rect 299944 205408 300264 216048
rect 306944 205408 307264 216048
rect 313944 205408 314264 216048
rect 320944 205408 321264 216048
rect 327944 205408 328264 216048
rect 334944 205408 335264 216048
rect 299944 149408 300264 160048
rect 306944 149408 307264 160048
rect 313944 149408 314264 160048
rect 320944 149408 321264 160048
rect 327944 149408 328264 160048
rect 334944 149408 335264 160048
rect 299944 93408 300264 104048
rect 306944 93408 307264 104048
rect 313944 93408 314264 104048
rect 320944 93408 321264 104048
rect 327944 93408 328264 104048
rect 334944 93408 335264 104048
rect 299944 156 300264 48048
rect 306944 156 307264 48048
rect 313944 156 314264 48048
rect 320944 156 321264 48048
rect 327944 156 328264 48048
rect 334944 156 335264 48048
rect 341944 156 342264 703780
rect 348944 156 349264 703780
rect 355944 653408 356264 703780
rect 362944 653408 363264 703780
rect 369944 653408 370264 703780
rect 376944 653408 377264 703780
rect 383944 653408 384264 703780
rect 390944 653408 391264 703780
rect 355944 597408 356264 608048
rect 362944 597408 363264 608048
rect 369944 597408 370264 608048
rect 376944 597408 377264 608048
rect 383944 597408 384264 608048
rect 390944 597408 391264 608048
rect 355944 541408 356264 552048
rect 362944 541408 363264 552048
rect 369944 541408 370264 552048
rect 376944 541408 377264 552048
rect 383944 541408 384264 552048
rect 390944 541408 391264 552048
rect 355944 485408 356264 496048
rect 362944 485408 363264 496048
rect 369944 485408 370264 496048
rect 376944 485408 377264 496048
rect 383944 485408 384264 496048
rect 390944 485408 391264 496048
rect 355944 429408 356264 440048
rect 362944 429408 363264 440048
rect 369944 429408 370264 440048
rect 376944 429408 377264 440048
rect 383944 429408 384264 440048
rect 390944 429408 391264 440048
rect 355944 373408 356264 384048
rect 362944 373408 363264 384048
rect 369944 373408 370264 384048
rect 376944 373408 377264 384048
rect 383944 373408 384264 384048
rect 390944 373408 391264 384048
rect 355944 317408 356264 328048
rect 362944 317408 363264 328048
rect 369944 317408 370264 328048
rect 376944 317408 377264 328048
rect 383944 317408 384264 328048
rect 390944 317408 391264 328048
rect 355944 261408 356264 272048
rect 362944 261408 363264 272048
rect 369944 261408 370264 272048
rect 376944 261408 377264 272048
rect 383944 261408 384264 272048
rect 390944 261408 391264 272048
rect 355944 205408 356264 216048
rect 362944 205408 363264 216048
rect 369944 205408 370264 216048
rect 376944 205408 377264 216048
rect 383944 205408 384264 216048
rect 390944 205408 391264 216048
rect 355944 149408 356264 160048
rect 362944 149408 363264 160048
rect 369944 149408 370264 160048
rect 376944 149408 377264 160048
rect 383944 149408 384264 160048
rect 390944 149408 391264 160048
rect 355944 93408 356264 104048
rect 362944 93408 363264 104048
rect 369944 93408 370264 104048
rect 376944 93408 377264 104048
rect 383944 93408 384264 104048
rect 390944 93408 391264 104048
rect 355944 156 356264 48048
rect 362944 156 363264 48048
rect 369944 156 370264 48048
rect 376944 156 377264 48048
rect 383944 156 384264 48048
rect 390944 156 391264 48048
rect 397944 156 398264 703780
rect 404944 156 405264 703780
rect 411944 653408 412264 703780
rect 418944 653408 419264 703780
rect 425944 653408 426264 703780
rect 432944 653408 433264 703780
rect 439944 653408 440264 703780
rect 446944 653408 447264 703780
rect 411944 597408 412264 608048
rect 418944 597408 419264 608048
rect 425944 597408 426264 608048
rect 432944 597408 433264 608048
rect 439944 597408 440264 608048
rect 446944 597408 447264 608048
rect 411944 541408 412264 552048
rect 418944 541408 419264 552048
rect 425944 541408 426264 552048
rect 432944 541408 433264 552048
rect 439944 541408 440264 552048
rect 446944 541408 447264 552048
rect 411944 485408 412264 496048
rect 418944 485408 419264 496048
rect 425944 485408 426264 496048
rect 432944 485408 433264 496048
rect 439944 485408 440264 496048
rect 446944 485408 447264 496048
rect 411944 429408 412264 440048
rect 418944 429408 419264 440048
rect 425944 429408 426264 440048
rect 432944 429408 433264 440048
rect 439944 429408 440264 440048
rect 446944 429408 447264 440048
rect 411944 373408 412264 384048
rect 418944 373408 419264 384048
rect 425944 373408 426264 384048
rect 432944 373408 433264 384048
rect 439944 373408 440264 384048
rect 446944 373408 447264 384048
rect 411944 317408 412264 328048
rect 418944 317408 419264 328048
rect 425944 317408 426264 328048
rect 432944 317408 433264 328048
rect 439944 317408 440264 328048
rect 446944 317408 447264 328048
rect 411944 261408 412264 272048
rect 418944 261408 419264 272048
rect 425944 261408 426264 272048
rect 432944 261408 433264 272048
rect 439944 261408 440264 272048
rect 446944 261408 447264 272048
rect 411944 205408 412264 216048
rect 418944 205408 419264 216048
rect 425944 205408 426264 216048
rect 432944 205408 433264 216048
rect 439944 205408 440264 216048
rect 446944 205408 447264 216048
rect 411944 149408 412264 160048
rect 418944 149408 419264 160048
rect 425944 149408 426264 160048
rect 432944 149408 433264 160048
rect 439944 149408 440264 160048
rect 446944 149408 447264 160048
rect 411944 93408 412264 104048
rect 418944 93408 419264 104048
rect 425944 93408 426264 104048
rect 432944 93408 433264 104048
rect 439944 93408 440264 104048
rect 446944 93408 447264 104048
rect 411944 156 412264 48048
rect 418944 156 419264 48048
rect 425944 156 426264 48048
rect 432944 156 433264 48048
rect 439944 156 440264 48048
rect 446944 156 447264 48048
rect 453944 156 454264 703780
rect 460944 156 461264 703780
rect 467944 653408 468264 703780
rect 474944 653408 475264 703780
rect 481944 653408 482264 703780
rect 488944 653408 489264 703780
rect 495944 653408 496264 703780
rect 502944 653408 503264 703780
rect 467944 597408 468264 608048
rect 474944 597408 475264 608048
rect 481944 597408 482264 608048
rect 488944 597408 489264 608048
rect 495944 597408 496264 608048
rect 502944 597408 503264 608048
rect 467944 541408 468264 552048
rect 474944 541408 475264 552048
rect 481944 541408 482264 552048
rect 488944 541408 489264 552048
rect 495944 541408 496264 552048
rect 502944 541408 503264 552048
rect 467944 485408 468264 496048
rect 474944 485408 475264 496048
rect 481944 485408 482264 496048
rect 488944 485408 489264 496048
rect 495944 485408 496264 496048
rect 502944 485408 503264 496048
rect 467944 429408 468264 440048
rect 474944 429408 475264 440048
rect 481944 429408 482264 440048
rect 488944 429408 489264 440048
rect 495944 429408 496264 440048
rect 502944 429408 503264 440048
rect 467944 373408 468264 384048
rect 474944 373408 475264 384048
rect 481944 373408 482264 384048
rect 488944 373408 489264 384048
rect 495944 373408 496264 384048
rect 502944 373408 503264 384048
rect 467944 317408 468264 328048
rect 474944 317408 475264 328048
rect 481944 317408 482264 328048
rect 488944 317408 489264 328048
rect 495944 317408 496264 328048
rect 502944 317408 503264 328048
rect 467944 261408 468264 272048
rect 474944 261408 475264 272048
rect 481944 261408 482264 272048
rect 488944 261408 489264 272048
rect 495944 261408 496264 272048
rect 502944 261408 503264 272048
rect 467944 205408 468264 216048
rect 474944 205408 475264 216048
rect 481944 205408 482264 216048
rect 488944 205408 489264 216048
rect 495944 205408 496264 216048
rect 502944 205408 503264 216048
rect 467944 149408 468264 160048
rect 474944 149408 475264 160048
rect 481944 149408 482264 160048
rect 488944 149408 489264 160048
rect 495944 149408 496264 160048
rect 502944 149408 503264 160048
rect 467944 93408 468264 104048
rect 474944 93408 475264 104048
rect 481944 93408 482264 104048
rect 488944 93408 489264 104048
rect 495944 93408 496264 104048
rect 502944 93408 503264 104048
rect 467944 156 468264 48048
rect 474944 156 475264 48048
rect 481944 156 482264 48048
rect 488944 156 489264 48048
rect 495944 156 496264 48048
rect 502944 156 503264 48048
rect 509944 156 510264 703780
rect 516944 156 517264 703780
rect 523944 653408 524264 703780
rect 530944 653408 531264 703780
rect 537944 653408 538264 703780
rect 544944 653408 545264 703780
rect 551944 653408 552264 703780
rect 558944 653408 559264 703780
rect 523944 597408 524264 608048
rect 530944 597408 531264 608048
rect 537944 597408 538264 608048
rect 544944 597408 545264 608048
rect 551944 597408 552264 608048
rect 558944 597408 559264 608048
rect 523944 541408 524264 552048
rect 530944 541408 531264 552048
rect 537944 541408 538264 552048
rect 544944 541408 545264 552048
rect 551944 541408 552264 552048
rect 558944 541408 559264 552048
rect 523944 485408 524264 496048
rect 530944 485408 531264 496048
rect 537944 485408 538264 496048
rect 544944 485408 545264 496048
rect 551944 485408 552264 496048
rect 558944 485408 559264 496048
rect 523944 429408 524264 440048
rect 530944 429408 531264 440048
rect 537944 429408 538264 440048
rect 544944 429408 545264 440048
rect 551944 429408 552264 440048
rect 558944 429408 559264 440048
rect 523944 373408 524264 384048
rect 530944 373408 531264 384048
rect 537944 373408 538264 384048
rect 544944 373408 545264 384048
rect 551944 373408 552264 384048
rect 558944 373408 559264 384048
rect 523944 317408 524264 328048
rect 530944 317408 531264 328048
rect 537944 317408 538264 328048
rect 544944 317408 545264 328048
rect 551944 317408 552264 328048
rect 558944 317408 559264 328048
rect 523944 261408 524264 272048
rect 530944 261408 531264 272048
rect 537944 261408 538264 272048
rect 544944 261408 545264 272048
rect 551944 261408 552264 272048
rect 558944 261408 559264 272048
rect 523944 205408 524264 216048
rect 530944 205408 531264 216048
rect 537944 205408 538264 216048
rect 544944 205408 545264 216048
rect 551944 205408 552264 216048
rect 558944 205408 559264 216048
rect 523944 149408 524264 160048
rect 530944 149408 531264 160048
rect 537944 149408 538264 160048
rect 544944 149408 545264 160048
rect 551944 149408 552264 160048
rect 558944 149408 559264 160048
rect 523944 93408 524264 104048
rect 530944 93408 531264 104048
rect 537944 93408 538264 104048
rect 544944 93408 545264 104048
rect 551944 93408 552264 104048
rect 558944 93408 559264 104048
rect 523944 156 524264 48048
rect 530944 156 531264 48048
rect 537944 156 538264 48048
rect 544944 156 545264 48048
rect 551944 156 552264 48048
rect 558944 156 559264 48048
rect 565944 156 566264 703780
rect 572944 156 573264 703780
rect 579944 156 580264 703780
rect 583860 816 584180 703120
rect 584520 156 584840 703780
<< obsm4 >>
rect 6499 2075 12864 655757
rect 13344 653328 19864 655757
rect 20344 653328 26864 655757
rect 27344 653328 33864 655757
rect 34344 653328 40864 655757
rect 41344 653328 47864 655757
rect 48344 653328 54864 655757
rect 55344 653328 61864 655757
rect 13344 608128 61864 653328
rect 13344 597328 19864 608128
rect 20344 597328 26864 608128
rect 27344 597328 33864 608128
rect 34344 597328 40864 608128
rect 41344 597328 47864 608128
rect 48344 597328 54864 608128
rect 55344 597328 61864 608128
rect 13344 552128 61864 597328
rect 13344 541328 19864 552128
rect 20344 541328 26864 552128
rect 27344 541328 33864 552128
rect 34344 541328 40864 552128
rect 41344 541328 47864 552128
rect 48344 541328 54864 552128
rect 55344 541328 61864 552128
rect 13344 496128 61864 541328
rect 13344 485328 19864 496128
rect 20344 485328 26864 496128
rect 27344 485328 33864 496128
rect 34344 485328 40864 496128
rect 41344 485328 47864 496128
rect 48344 485328 54864 496128
rect 55344 485328 61864 496128
rect 13344 440128 61864 485328
rect 13344 429328 19864 440128
rect 20344 429328 26864 440128
rect 27344 429328 33864 440128
rect 34344 429328 40864 440128
rect 41344 429328 47864 440128
rect 48344 429328 54864 440128
rect 55344 429328 61864 440128
rect 13344 384128 61864 429328
rect 13344 373328 19864 384128
rect 20344 373328 26864 384128
rect 27344 373328 33864 384128
rect 34344 373328 40864 384128
rect 41344 373328 47864 384128
rect 48344 373328 54864 384128
rect 55344 373328 61864 384128
rect 13344 328128 61864 373328
rect 13344 317328 19864 328128
rect 20344 317328 26864 328128
rect 27344 317328 33864 328128
rect 34344 317328 40864 328128
rect 41344 317328 47864 328128
rect 48344 317328 54864 328128
rect 55344 317328 61864 328128
rect 13344 272128 61864 317328
rect 13344 261328 19864 272128
rect 20344 261328 26864 272128
rect 27344 261328 33864 272128
rect 34344 261328 40864 272128
rect 41344 261328 47864 272128
rect 48344 261328 54864 272128
rect 55344 261328 61864 272128
rect 13344 216128 61864 261328
rect 13344 205328 19864 216128
rect 20344 205328 26864 216128
rect 27344 205328 33864 216128
rect 34344 205328 40864 216128
rect 41344 205328 47864 216128
rect 48344 205328 54864 216128
rect 55344 205328 61864 216128
rect 13344 160128 61864 205328
rect 13344 149328 19864 160128
rect 20344 149328 26864 160128
rect 27344 149328 33864 160128
rect 34344 149328 40864 160128
rect 41344 149328 47864 160128
rect 48344 149328 54864 160128
rect 55344 149328 61864 160128
rect 13344 104128 61864 149328
rect 13344 93328 19864 104128
rect 20344 93328 26864 104128
rect 27344 93328 33864 104128
rect 34344 93328 40864 104128
rect 41344 93328 47864 104128
rect 48344 93328 54864 104128
rect 55344 93328 61864 104128
rect 13344 48128 61864 93328
rect 13344 2075 19864 48128
rect 20344 2075 26864 48128
rect 27344 2075 33864 48128
rect 34344 2075 40864 48128
rect 41344 2075 47864 48128
rect 48344 2075 54864 48128
rect 55344 2075 61864 48128
rect 62344 2075 68864 655757
rect 69344 653328 75864 655757
rect 76344 653328 82864 655757
rect 83344 653328 89864 655757
rect 90344 653328 96864 655757
rect 97344 653328 103864 655757
rect 104344 653328 110864 655757
rect 111344 653328 117864 655757
rect 69344 608128 117864 653328
rect 69344 597328 75864 608128
rect 76344 597328 82864 608128
rect 83344 597328 89864 608128
rect 90344 597328 96864 608128
rect 97344 597328 103864 608128
rect 104344 597328 110864 608128
rect 111344 597328 117864 608128
rect 69344 552128 117864 597328
rect 69344 541328 75864 552128
rect 76344 541328 82864 552128
rect 83344 541328 89864 552128
rect 90344 541328 96864 552128
rect 97344 541328 103864 552128
rect 104344 541328 110864 552128
rect 111344 541328 117864 552128
rect 69344 496128 117864 541328
rect 69344 485328 75864 496128
rect 76344 485328 82864 496128
rect 83344 485328 89864 496128
rect 90344 485328 96864 496128
rect 97344 485328 103864 496128
rect 104344 485328 110864 496128
rect 111344 485328 117864 496128
rect 69344 440128 117864 485328
rect 69344 429328 75864 440128
rect 76344 429328 82864 440128
rect 83344 429328 89864 440128
rect 90344 429328 96864 440128
rect 97344 429328 103864 440128
rect 104344 429328 110864 440128
rect 111344 429328 117864 440128
rect 69344 384128 117864 429328
rect 69344 373328 75864 384128
rect 76344 373328 82864 384128
rect 83344 373328 89864 384128
rect 90344 373328 96864 384128
rect 97344 373328 103864 384128
rect 104344 373328 110864 384128
rect 111344 373328 117864 384128
rect 69344 328128 117864 373328
rect 69344 317328 75864 328128
rect 76344 317328 82864 328128
rect 83344 317328 89864 328128
rect 90344 317328 96864 328128
rect 97344 317328 103864 328128
rect 104344 317328 110864 328128
rect 111344 317328 117864 328128
rect 69344 272128 117864 317328
rect 69344 261328 75864 272128
rect 76344 261328 82864 272128
rect 83344 261328 89864 272128
rect 90344 261328 96864 272128
rect 97344 261328 103864 272128
rect 104344 261328 110864 272128
rect 111344 261328 117864 272128
rect 69344 216128 117864 261328
rect 69344 205328 75864 216128
rect 76344 205328 82864 216128
rect 83344 205328 89864 216128
rect 90344 205328 96864 216128
rect 97344 205328 103864 216128
rect 104344 205328 110864 216128
rect 111344 205328 117864 216128
rect 69344 160128 117864 205328
rect 69344 149328 75864 160128
rect 76344 149328 82864 160128
rect 83344 149328 89864 160128
rect 90344 149328 96864 160128
rect 97344 149328 103864 160128
rect 104344 149328 110864 160128
rect 111344 149328 117864 160128
rect 69344 104128 117864 149328
rect 69344 93328 75864 104128
rect 76344 93328 82864 104128
rect 83344 93328 89864 104128
rect 90344 93328 96864 104128
rect 97344 93328 103864 104128
rect 104344 93328 110864 104128
rect 111344 93328 117864 104128
rect 69344 48128 117864 93328
rect 69344 2075 75864 48128
rect 76344 2075 82864 48128
rect 83344 2075 89864 48128
rect 90344 2075 96864 48128
rect 97344 2075 103864 48128
rect 104344 2075 110864 48128
rect 111344 2075 117864 48128
rect 118344 2075 124864 655757
rect 125344 653328 131864 655757
rect 132344 653328 138864 655757
rect 139344 653328 145864 655757
rect 146344 653328 152864 655757
rect 153344 653328 159864 655757
rect 160344 653328 166864 655757
rect 167344 653328 173864 655757
rect 125344 608128 173864 653328
rect 125344 597328 131864 608128
rect 132344 597328 138864 608128
rect 139344 597328 145864 608128
rect 146344 597328 152864 608128
rect 153344 597328 159864 608128
rect 160344 597328 166864 608128
rect 167344 597328 173864 608128
rect 125344 552128 173864 597328
rect 125344 541328 131864 552128
rect 132344 541328 138864 552128
rect 139344 541328 145864 552128
rect 146344 541328 152864 552128
rect 153344 541328 159864 552128
rect 160344 541328 166864 552128
rect 167344 541328 173864 552128
rect 125344 496128 173864 541328
rect 125344 485328 131864 496128
rect 132344 485328 138864 496128
rect 139344 485328 145864 496128
rect 146344 485328 152864 496128
rect 153344 485328 159864 496128
rect 160344 485328 166864 496128
rect 167344 485328 173864 496128
rect 125344 440128 173864 485328
rect 125344 429328 131864 440128
rect 132344 429328 138864 440128
rect 139344 429328 145864 440128
rect 146344 429328 152864 440128
rect 153344 429328 159864 440128
rect 160344 429328 166864 440128
rect 167344 429328 173864 440128
rect 125344 384128 173864 429328
rect 125344 373328 131864 384128
rect 132344 373328 138864 384128
rect 139344 373328 145864 384128
rect 146344 373328 152864 384128
rect 153344 373328 159864 384128
rect 160344 373328 166864 384128
rect 167344 373328 173864 384128
rect 125344 328128 173864 373328
rect 125344 317328 131864 328128
rect 132344 317328 138864 328128
rect 139344 317328 145864 328128
rect 146344 317328 152864 328128
rect 153344 317328 159864 328128
rect 160344 317328 166864 328128
rect 167344 317328 173864 328128
rect 125344 272128 173864 317328
rect 125344 261328 131864 272128
rect 132344 261328 138864 272128
rect 139344 261328 145864 272128
rect 146344 261328 152864 272128
rect 153344 261328 159864 272128
rect 160344 261328 166864 272128
rect 167344 261328 173864 272128
rect 125344 216128 173864 261328
rect 125344 205328 131864 216128
rect 132344 205328 138864 216128
rect 139344 205328 145864 216128
rect 146344 205328 152864 216128
rect 153344 205328 159864 216128
rect 160344 205328 166864 216128
rect 167344 205328 173864 216128
rect 125344 160128 173864 205328
rect 125344 149328 131864 160128
rect 132344 149328 138864 160128
rect 139344 149328 145864 160128
rect 146344 149328 152864 160128
rect 153344 149328 159864 160128
rect 160344 149328 166864 160128
rect 167344 149328 173864 160128
rect 125344 104128 173864 149328
rect 125344 93328 131864 104128
rect 132344 93328 138864 104128
rect 139344 93328 145864 104128
rect 146344 93328 152864 104128
rect 153344 93328 159864 104128
rect 160344 93328 166864 104128
rect 167344 93328 173864 104128
rect 125344 48128 173864 93328
rect 125344 2075 131864 48128
rect 132344 2075 138864 48128
rect 139344 2075 145864 48128
rect 146344 2075 152864 48128
rect 153344 2075 159864 48128
rect 160344 2075 166864 48128
rect 167344 2075 173864 48128
rect 174344 2075 180864 655757
rect 181344 653328 187864 655757
rect 188344 653328 194864 655757
rect 195344 653328 201864 655757
rect 202344 653328 208864 655757
rect 209344 653328 215864 655757
rect 216344 653328 222864 655757
rect 223344 653328 229864 655757
rect 181344 608128 229864 653328
rect 181344 597328 187864 608128
rect 188344 597328 194864 608128
rect 195344 597328 201864 608128
rect 202344 597328 208864 608128
rect 209344 597328 215864 608128
rect 216344 597328 222864 608128
rect 223344 597328 229864 608128
rect 181344 552128 229864 597328
rect 181344 541328 187864 552128
rect 188344 541328 194864 552128
rect 195344 541328 201864 552128
rect 202344 541328 208864 552128
rect 209344 541328 215864 552128
rect 216344 541328 222864 552128
rect 223344 541328 229864 552128
rect 181344 496128 229864 541328
rect 181344 485328 187864 496128
rect 188344 485328 194864 496128
rect 195344 485328 201864 496128
rect 202344 485328 208864 496128
rect 209344 485328 215864 496128
rect 216344 485328 222864 496128
rect 223344 485328 229864 496128
rect 181344 440128 229864 485328
rect 181344 429328 187864 440128
rect 188344 429328 194864 440128
rect 195344 429328 201864 440128
rect 202344 429328 208864 440128
rect 209344 429328 215864 440128
rect 216344 429328 222864 440128
rect 223344 429328 229864 440128
rect 181344 384128 229864 429328
rect 181344 373328 187864 384128
rect 188344 373328 194864 384128
rect 195344 373328 201864 384128
rect 202344 373328 208864 384128
rect 209344 373328 215864 384128
rect 216344 373328 222864 384128
rect 223344 373328 229864 384128
rect 181344 328128 229864 373328
rect 181344 317328 187864 328128
rect 188344 317328 194864 328128
rect 195344 317328 201864 328128
rect 202344 317328 208864 328128
rect 209344 317328 215864 328128
rect 216344 317328 222864 328128
rect 223344 317328 229864 328128
rect 181344 272128 229864 317328
rect 181344 261328 187864 272128
rect 188344 261328 194864 272128
rect 195344 261328 201864 272128
rect 202344 261328 208864 272128
rect 209344 261328 215864 272128
rect 216344 261328 222864 272128
rect 223344 261328 229864 272128
rect 181344 216128 229864 261328
rect 181344 205328 187864 216128
rect 188344 205328 194864 216128
rect 195344 205328 201864 216128
rect 202344 205328 208864 216128
rect 209344 205328 215864 216128
rect 216344 205328 222864 216128
rect 223344 205328 229864 216128
rect 181344 160128 229864 205328
rect 181344 149328 187864 160128
rect 188344 149328 194864 160128
rect 195344 149328 201864 160128
rect 202344 149328 208864 160128
rect 209344 149328 215864 160128
rect 216344 149328 222864 160128
rect 223344 149328 229864 160128
rect 181344 104128 229864 149328
rect 181344 93328 187864 104128
rect 188344 93328 194864 104128
rect 195344 93328 201864 104128
rect 202344 93328 208864 104128
rect 209344 93328 215864 104128
rect 216344 93328 222864 104128
rect 223344 93328 229864 104128
rect 181344 48128 229864 93328
rect 181344 2075 187864 48128
rect 188344 2075 194864 48128
rect 195344 2075 201864 48128
rect 202344 2075 208864 48128
rect 209344 2075 215864 48128
rect 216344 2075 222864 48128
rect 223344 2075 229864 48128
rect 230344 2075 236864 655757
rect 237344 653328 243864 655757
rect 244344 653328 250864 655757
rect 251344 653328 257864 655757
rect 258344 653328 264864 655757
rect 265344 653328 271864 655757
rect 272344 653328 278864 655757
rect 279344 653328 285864 655757
rect 237344 608128 285864 653328
rect 237344 597328 243864 608128
rect 244344 597328 250864 608128
rect 251344 597328 257864 608128
rect 258344 597328 264864 608128
rect 265344 597328 271864 608128
rect 272344 597328 278864 608128
rect 279344 597328 285864 608128
rect 237344 552128 285864 597328
rect 237344 541328 243864 552128
rect 244344 541328 250864 552128
rect 251344 541328 257864 552128
rect 258344 541328 264864 552128
rect 265344 541328 271864 552128
rect 272344 541328 278864 552128
rect 279344 541328 285864 552128
rect 237344 496128 285864 541328
rect 237344 485328 243864 496128
rect 244344 485328 250864 496128
rect 251344 485328 257864 496128
rect 258344 485328 264864 496128
rect 265344 485328 271864 496128
rect 272344 485328 278864 496128
rect 279344 485328 285864 496128
rect 237344 440128 285864 485328
rect 237344 429328 243864 440128
rect 244344 429328 250864 440128
rect 251344 429328 257864 440128
rect 258344 429328 264864 440128
rect 265344 429328 271864 440128
rect 272344 429328 278864 440128
rect 279344 429328 285864 440128
rect 237344 384128 285864 429328
rect 237344 373328 243864 384128
rect 244344 373328 250864 384128
rect 251344 373328 257864 384128
rect 258344 373328 264864 384128
rect 265344 373328 271864 384128
rect 272344 373328 278864 384128
rect 279344 373328 285864 384128
rect 237344 328128 285864 373328
rect 237344 317328 243864 328128
rect 244344 317328 250864 328128
rect 251344 317328 257864 328128
rect 258344 317328 264864 328128
rect 265344 317328 271864 328128
rect 272344 317328 278864 328128
rect 279344 317328 285864 328128
rect 237344 272128 285864 317328
rect 237344 261328 243864 272128
rect 244344 261328 250864 272128
rect 251344 261328 257864 272128
rect 258344 261328 264864 272128
rect 265344 261328 271864 272128
rect 272344 261328 278864 272128
rect 279344 261328 285864 272128
rect 237344 216128 285864 261328
rect 237344 205328 243864 216128
rect 244344 205328 250864 216128
rect 251344 205328 257864 216128
rect 258344 205328 264864 216128
rect 265344 205328 271864 216128
rect 272344 205328 278864 216128
rect 279344 205328 285864 216128
rect 237344 160128 285864 205328
rect 237344 149328 243864 160128
rect 244344 149328 250864 160128
rect 251344 149328 257864 160128
rect 258344 149328 264864 160128
rect 265344 149328 271864 160128
rect 272344 149328 278864 160128
rect 279344 149328 285864 160128
rect 237344 104128 285864 149328
rect 237344 93328 243864 104128
rect 244344 93328 250864 104128
rect 251344 93328 257864 104128
rect 258344 93328 264864 104128
rect 265344 93328 271864 104128
rect 272344 93328 278864 104128
rect 279344 93328 285864 104128
rect 237344 48128 285864 93328
rect 237344 2075 243864 48128
rect 244344 2075 250864 48128
rect 251344 2075 257864 48128
rect 258344 2075 264864 48128
rect 265344 2075 271864 48128
rect 272344 2075 278864 48128
rect 279344 2075 285864 48128
rect 286344 2075 292864 655757
rect 293344 653328 299864 655757
rect 300344 653328 306864 655757
rect 307344 653328 313864 655757
rect 314344 653328 320864 655757
rect 321344 653328 327864 655757
rect 328344 653328 334864 655757
rect 335344 653328 341864 655757
rect 293344 608128 341864 653328
rect 293344 597328 299864 608128
rect 300344 597328 306864 608128
rect 307344 597328 313864 608128
rect 314344 597328 320864 608128
rect 321344 597328 327864 608128
rect 328344 597328 334864 608128
rect 335344 597328 341864 608128
rect 293344 552128 341864 597328
rect 293344 541328 299864 552128
rect 300344 541328 306864 552128
rect 307344 541328 313864 552128
rect 314344 541328 320864 552128
rect 321344 541328 327864 552128
rect 328344 541328 334864 552128
rect 335344 541328 341864 552128
rect 293344 496128 341864 541328
rect 293344 485328 299864 496128
rect 300344 485328 306864 496128
rect 307344 485328 313864 496128
rect 314344 485328 320864 496128
rect 321344 485328 327864 496128
rect 328344 485328 334864 496128
rect 335344 485328 341864 496128
rect 293344 440128 341864 485328
rect 293344 429328 299864 440128
rect 300344 429328 306864 440128
rect 307344 429328 313864 440128
rect 314344 429328 320864 440128
rect 321344 429328 327864 440128
rect 328344 429328 334864 440128
rect 335344 429328 341864 440128
rect 293344 384128 341864 429328
rect 293344 373328 299864 384128
rect 300344 373328 306864 384128
rect 307344 373328 313864 384128
rect 314344 373328 320864 384128
rect 321344 373328 327864 384128
rect 328344 373328 334864 384128
rect 335344 373328 341864 384128
rect 293344 328128 341864 373328
rect 293344 317328 299864 328128
rect 300344 317328 306864 328128
rect 307344 317328 313864 328128
rect 314344 317328 320864 328128
rect 321344 317328 327864 328128
rect 328344 317328 334864 328128
rect 335344 317328 341864 328128
rect 293344 272128 341864 317328
rect 293344 261328 299864 272128
rect 300344 261328 306864 272128
rect 307344 261328 313864 272128
rect 314344 261328 320864 272128
rect 321344 261328 327864 272128
rect 328344 261328 334864 272128
rect 335344 261328 341864 272128
rect 293344 216128 341864 261328
rect 293344 205328 299864 216128
rect 300344 205328 306864 216128
rect 307344 205328 313864 216128
rect 314344 205328 320864 216128
rect 321344 205328 327864 216128
rect 328344 205328 334864 216128
rect 335344 205328 341864 216128
rect 293344 160128 341864 205328
rect 293344 149328 299864 160128
rect 300344 149328 306864 160128
rect 307344 149328 313864 160128
rect 314344 149328 320864 160128
rect 321344 149328 327864 160128
rect 328344 149328 334864 160128
rect 335344 149328 341864 160128
rect 293344 104128 341864 149328
rect 293344 93328 299864 104128
rect 300344 93328 306864 104128
rect 307344 93328 313864 104128
rect 314344 93328 320864 104128
rect 321344 93328 327864 104128
rect 328344 93328 334864 104128
rect 335344 93328 341864 104128
rect 293344 48128 341864 93328
rect 293344 2075 299864 48128
rect 300344 2075 306864 48128
rect 307344 2075 313864 48128
rect 314344 2075 320864 48128
rect 321344 2075 327864 48128
rect 328344 2075 334864 48128
rect 335344 2075 341864 48128
rect 342344 2075 348864 655757
rect 349344 653328 355864 655757
rect 356344 653328 362864 655757
rect 363344 653328 369864 655757
rect 370344 653328 376864 655757
rect 377344 653328 383864 655757
rect 384344 653328 390864 655757
rect 391344 653328 397864 655757
rect 349344 608128 397864 653328
rect 349344 597328 355864 608128
rect 356344 597328 362864 608128
rect 363344 597328 369864 608128
rect 370344 597328 376864 608128
rect 377344 597328 383864 608128
rect 384344 597328 390864 608128
rect 391344 597328 397864 608128
rect 349344 552128 397864 597328
rect 349344 541328 355864 552128
rect 356344 541328 362864 552128
rect 363344 541328 369864 552128
rect 370344 541328 376864 552128
rect 377344 541328 383864 552128
rect 384344 541328 390864 552128
rect 391344 541328 397864 552128
rect 349344 496128 397864 541328
rect 349344 485328 355864 496128
rect 356344 485328 362864 496128
rect 363344 485328 369864 496128
rect 370344 485328 376864 496128
rect 377344 485328 383864 496128
rect 384344 485328 390864 496128
rect 391344 485328 397864 496128
rect 349344 440128 397864 485328
rect 349344 429328 355864 440128
rect 356344 429328 362864 440128
rect 363344 429328 369864 440128
rect 370344 429328 376864 440128
rect 377344 429328 383864 440128
rect 384344 429328 390864 440128
rect 391344 429328 397864 440128
rect 349344 384128 397864 429328
rect 349344 373328 355864 384128
rect 356344 373328 362864 384128
rect 363344 373328 369864 384128
rect 370344 373328 376864 384128
rect 377344 373328 383864 384128
rect 384344 373328 390864 384128
rect 391344 373328 397864 384128
rect 349344 328128 397864 373328
rect 349344 317328 355864 328128
rect 356344 317328 362864 328128
rect 363344 317328 369864 328128
rect 370344 317328 376864 328128
rect 377344 317328 383864 328128
rect 384344 317328 390864 328128
rect 391344 317328 397864 328128
rect 349344 272128 397864 317328
rect 349344 261328 355864 272128
rect 356344 261328 362864 272128
rect 363344 261328 369864 272128
rect 370344 261328 376864 272128
rect 377344 261328 383864 272128
rect 384344 261328 390864 272128
rect 391344 261328 397864 272128
rect 349344 216128 397864 261328
rect 349344 205328 355864 216128
rect 356344 205328 362864 216128
rect 363344 205328 369864 216128
rect 370344 205328 376864 216128
rect 377344 205328 383864 216128
rect 384344 205328 390864 216128
rect 391344 205328 397864 216128
rect 349344 160128 397864 205328
rect 349344 149328 355864 160128
rect 356344 149328 362864 160128
rect 363344 149328 369864 160128
rect 370344 149328 376864 160128
rect 377344 149328 383864 160128
rect 384344 149328 390864 160128
rect 391344 149328 397864 160128
rect 349344 104128 397864 149328
rect 349344 93328 355864 104128
rect 356344 93328 362864 104128
rect 363344 93328 369864 104128
rect 370344 93328 376864 104128
rect 377344 93328 383864 104128
rect 384344 93328 390864 104128
rect 391344 93328 397864 104128
rect 349344 48128 397864 93328
rect 349344 2075 355864 48128
rect 356344 2075 362864 48128
rect 363344 2075 369864 48128
rect 370344 2075 376864 48128
rect 377344 2075 383864 48128
rect 384344 2075 390864 48128
rect 391344 2075 397864 48128
rect 398344 2075 404864 655757
rect 405344 653328 411864 655757
rect 412344 653328 418864 655757
rect 419344 653328 425864 655757
rect 426344 653328 432864 655757
rect 433344 653328 439864 655757
rect 440344 653328 446864 655757
rect 447344 653328 453864 655757
rect 405344 608128 453864 653328
rect 405344 597328 411864 608128
rect 412344 597328 418864 608128
rect 419344 597328 425864 608128
rect 426344 597328 432864 608128
rect 433344 597328 439864 608128
rect 440344 597328 446864 608128
rect 447344 597328 453864 608128
rect 405344 552128 453864 597328
rect 405344 541328 411864 552128
rect 412344 541328 418864 552128
rect 419344 541328 425864 552128
rect 426344 541328 432864 552128
rect 433344 541328 439864 552128
rect 440344 541328 446864 552128
rect 447344 541328 453864 552128
rect 405344 496128 453864 541328
rect 405344 485328 411864 496128
rect 412344 485328 418864 496128
rect 419344 485328 425864 496128
rect 426344 485328 432864 496128
rect 433344 485328 439864 496128
rect 440344 485328 446864 496128
rect 447344 485328 453864 496128
rect 405344 440128 453864 485328
rect 405344 429328 411864 440128
rect 412344 429328 418864 440128
rect 419344 429328 425864 440128
rect 426344 429328 432864 440128
rect 433344 429328 439864 440128
rect 440344 429328 446864 440128
rect 447344 429328 453864 440128
rect 405344 384128 453864 429328
rect 405344 373328 411864 384128
rect 412344 373328 418864 384128
rect 419344 373328 425864 384128
rect 426344 373328 432864 384128
rect 433344 373328 439864 384128
rect 440344 373328 446864 384128
rect 447344 373328 453864 384128
rect 405344 328128 453864 373328
rect 405344 317328 411864 328128
rect 412344 317328 418864 328128
rect 419344 317328 425864 328128
rect 426344 317328 432864 328128
rect 433344 317328 439864 328128
rect 440344 317328 446864 328128
rect 447344 317328 453864 328128
rect 405344 272128 453864 317328
rect 405344 261328 411864 272128
rect 412344 261328 418864 272128
rect 419344 261328 425864 272128
rect 426344 261328 432864 272128
rect 433344 261328 439864 272128
rect 440344 261328 446864 272128
rect 447344 261328 453864 272128
rect 405344 216128 453864 261328
rect 405344 205328 411864 216128
rect 412344 205328 418864 216128
rect 419344 205328 425864 216128
rect 426344 205328 432864 216128
rect 433344 205328 439864 216128
rect 440344 205328 446864 216128
rect 447344 205328 453864 216128
rect 405344 160128 453864 205328
rect 405344 149328 411864 160128
rect 412344 149328 418864 160128
rect 419344 149328 425864 160128
rect 426344 149328 432864 160128
rect 433344 149328 439864 160128
rect 440344 149328 446864 160128
rect 447344 149328 453864 160128
rect 405344 104128 453864 149328
rect 405344 93328 411864 104128
rect 412344 93328 418864 104128
rect 419344 93328 425864 104128
rect 426344 93328 432864 104128
rect 433344 93328 439864 104128
rect 440344 93328 446864 104128
rect 447344 93328 453864 104128
rect 405344 48128 453864 93328
rect 405344 2075 411864 48128
rect 412344 2075 418864 48128
rect 419344 2075 425864 48128
rect 426344 2075 432864 48128
rect 433344 2075 439864 48128
rect 440344 2075 446864 48128
rect 447344 2075 453864 48128
rect 454344 2075 460864 655757
rect 461344 653328 467864 655757
rect 468344 653328 474864 655757
rect 475344 653328 481864 655757
rect 482344 653328 488864 655757
rect 489344 653328 495864 655757
rect 496344 653328 502864 655757
rect 503344 653328 509864 655757
rect 461344 608128 509864 653328
rect 461344 597328 467864 608128
rect 468344 597328 474864 608128
rect 475344 597328 481864 608128
rect 482344 597328 488864 608128
rect 489344 597328 495864 608128
rect 496344 597328 502864 608128
rect 503344 597328 509864 608128
rect 461344 552128 509864 597328
rect 461344 541328 467864 552128
rect 468344 541328 474864 552128
rect 475344 541328 481864 552128
rect 482344 541328 488864 552128
rect 489344 541328 495864 552128
rect 496344 541328 502864 552128
rect 503344 541328 509864 552128
rect 461344 496128 509864 541328
rect 461344 485328 467864 496128
rect 468344 485328 474864 496128
rect 475344 485328 481864 496128
rect 482344 485328 488864 496128
rect 489344 485328 495864 496128
rect 496344 485328 502864 496128
rect 503344 485328 509864 496128
rect 461344 440128 509864 485328
rect 461344 429328 467864 440128
rect 468344 429328 474864 440128
rect 475344 429328 481864 440128
rect 482344 429328 488864 440128
rect 489344 429328 495864 440128
rect 496344 429328 502864 440128
rect 503344 429328 509864 440128
rect 461344 384128 509864 429328
rect 461344 373328 467864 384128
rect 468344 373328 474864 384128
rect 475344 373328 481864 384128
rect 482344 373328 488864 384128
rect 489344 373328 495864 384128
rect 496344 373328 502864 384128
rect 503344 373328 509864 384128
rect 461344 328128 509864 373328
rect 461344 317328 467864 328128
rect 468344 317328 474864 328128
rect 475344 317328 481864 328128
rect 482344 317328 488864 328128
rect 489344 317328 495864 328128
rect 496344 317328 502864 328128
rect 503344 317328 509864 328128
rect 461344 272128 509864 317328
rect 461344 261328 467864 272128
rect 468344 261328 474864 272128
rect 475344 261328 481864 272128
rect 482344 261328 488864 272128
rect 489344 261328 495864 272128
rect 496344 261328 502864 272128
rect 503344 261328 509864 272128
rect 461344 216128 509864 261328
rect 461344 205328 467864 216128
rect 468344 205328 474864 216128
rect 475344 205328 481864 216128
rect 482344 205328 488864 216128
rect 489344 205328 495864 216128
rect 496344 205328 502864 216128
rect 503344 205328 509864 216128
rect 461344 160128 509864 205328
rect 461344 149328 467864 160128
rect 468344 149328 474864 160128
rect 475344 149328 481864 160128
rect 482344 149328 488864 160128
rect 489344 149328 495864 160128
rect 496344 149328 502864 160128
rect 503344 149328 509864 160128
rect 461344 104128 509864 149328
rect 461344 93328 467864 104128
rect 468344 93328 474864 104128
rect 475344 93328 481864 104128
rect 482344 93328 488864 104128
rect 489344 93328 495864 104128
rect 496344 93328 502864 104128
rect 503344 93328 509864 104128
rect 461344 48128 509864 93328
rect 461344 2075 467864 48128
rect 468344 2075 474864 48128
rect 475344 2075 481864 48128
rect 482344 2075 488864 48128
rect 489344 2075 495864 48128
rect 496344 2075 502864 48128
rect 503344 2075 509864 48128
rect 510344 2075 516864 655757
rect 517344 653328 523864 655757
rect 524344 653328 530864 655757
rect 531344 653328 537864 655757
rect 538344 653328 544864 655757
rect 545344 653328 551864 655757
rect 552344 653328 558864 655757
rect 559344 653328 565864 655757
rect 517344 608128 565864 653328
rect 517344 597328 523864 608128
rect 524344 597328 530864 608128
rect 531344 597328 537864 608128
rect 538344 597328 544864 608128
rect 545344 597328 551864 608128
rect 552344 597328 558864 608128
rect 559344 597328 565864 608128
rect 517344 552128 565864 597328
rect 517344 541328 523864 552128
rect 524344 541328 530864 552128
rect 531344 541328 537864 552128
rect 538344 541328 544864 552128
rect 545344 541328 551864 552128
rect 552344 541328 558864 552128
rect 559344 541328 565864 552128
rect 517344 496128 565864 541328
rect 517344 485328 523864 496128
rect 524344 485328 530864 496128
rect 531344 485328 537864 496128
rect 538344 485328 544864 496128
rect 545344 485328 551864 496128
rect 552344 485328 558864 496128
rect 559344 485328 565864 496128
rect 517344 440128 565864 485328
rect 517344 429328 523864 440128
rect 524344 429328 530864 440128
rect 531344 429328 537864 440128
rect 538344 429328 544864 440128
rect 545344 429328 551864 440128
rect 552344 429328 558864 440128
rect 559344 429328 565864 440128
rect 517344 384128 565864 429328
rect 517344 373328 523864 384128
rect 524344 373328 530864 384128
rect 531344 373328 537864 384128
rect 538344 373328 544864 384128
rect 545344 373328 551864 384128
rect 552344 373328 558864 384128
rect 559344 373328 565864 384128
rect 517344 328128 565864 373328
rect 517344 317328 523864 328128
rect 524344 317328 530864 328128
rect 531344 317328 537864 328128
rect 538344 317328 544864 328128
rect 545344 317328 551864 328128
rect 552344 317328 558864 328128
rect 559344 317328 565864 328128
rect 517344 272128 565864 317328
rect 517344 261328 523864 272128
rect 524344 261328 530864 272128
rect 531344 261328 537864 272128
rect 538344 261328 544864 272128
rect 545344 261328 551864 272128
rect 552344 261328 558864 272128
rect 559344 261328 565864 272128
rect 517344 216128 565864 261328
rect 517344 205328 523864 216128
rect 524344 205328 530864 216128
rect 531344 205328 537864 216128
rect 538344 205328 544864 216128
rect 545344 205328 551864 216128
rect 552344 205328 558864 216128
rect 559344 205328 565864 216128
rect 517344 160128 565864 205328
rect 517344 149328 523864 160128
rect 524344 149328 530864 160128
rect 531344 149328 537864 160128
rect 538344 149328 544864 160128
rect 545344 149328 551864 160128
rect 552344 149328 558864 160128
rect 559344 149328 565864 160128
rect 517344 104128 565864 149328
rect 517344 93328 523864 104128
rect 524344 93328 530864 104128
rect 531344 93328 537864 104128
rect 538344 93328 544864 104128
rect 545344 93328 551864 104128
rect 552344 93328 558864 104128
rect 559344 93328 565864 104128
rect 517344 48128 565864 93328
rect 517344 2075 523864 48128
rect 524344 2075 530864 48128
rect 531344 2075 537864 48128
rect 538344 2075 544864 48128
rect 545344 2075 551864 48128
rect 552344 2075 558864 48128
rect 559344 2075 565864 48128
rect 566344 2075 572864 655757
rect 573344 2075 573837 655757
<< metal5 >>
rect -916 703460 584840 703780
rect -256 702800 584180 703120
rect -916 697968 584840 698288
rect -916 690968 584840 691288
rect -916 683968 584840 684288
rect -916 676968 584840 677288
rect -916 669968 584840 670288
rect -916 662968 584840 663288
rect -916 655968 584840 656288
rect -916 648968 584840 649288
rect -916 641968 584840 642288
rect -916 634968 584840 635288
rect -916 627968 584840 628288
rect -916 620968 584840 621288
rect -916 613968 584840 614288
rect -916 606968 584840 607288
rect -916 599968 584840 600288
rect -916 592968 584840 593288
rect -916 585968 584840 586288
rect -916 578968 584840 579288
rect -916 571968 584840 572288
rect -916 564968 584840 565288
rect -916 557968 584840 558288
rect -916 550968 584840 551288
rect -916 543968 584840 544288
rect -916 536968 584840 537288
rect -916 529968 584840 530288
rect -916 522968 584840 523288
rect -916 515968 584840 516288
rect -916 508968 584840 509288
rect -916 501968 584840 502288
rect -916 494968 584840 495288
rect -916 487968 584840 488288
rect -916 480968 584840 481288
rect -916 473968 584840 474288
rect -916 466968 584840 467288
rect -916 459968 584840 460288
rect -916 452968 584840 453288
rect -916 445968 584840 446288
rect -916 438968 584840 439288
rect -916 431968 584840 432288
rect -916 424968 584840 425288
rect -916 417968 584840 418288
rect -916 410968 584840 411288
rect -916 403968 584840 404288
rect -916 396968 584840 397288
rect -916 389968 584840 390288
rect -916 382968 584840 383288
rect -916 375968 584840 376288
rect -916 368968 584840 369288
rect -916 361968 584840 362288
rect -916 354968 584840 355288
rect -916 347968 584840 348288
rect -916 340968 584840 341288
rect -916 333968 584840 334288
rect -916 326968 584840 327288
rect -916 319968 584840 320288
rect -916 312968 584840 313288
rect -916 305968 584840 306288
rect -916 298968 584840 299288
rect -916 291968 584840 292288
rect -916 284968 584840 285288
rect -916 277968 584840 278288
rect -916 270968 584840 271288
rect -916 263968 584840 264288
rect -916 256968 584840 257288
rect -916 249968 584840 250288
rect -916 242968 584840 243288
rect -916 235968 584840 236288
rect -916 228968 584840 229288
rect -916 221968 584840 222288
rect -916 214968 584840 215288
rect -916 207968 584840 208288
rect -916 200968 584840 201288
rect -916 193968 584840 194288
rect -916 186968 584840 187288
rect -916 179968 584840 180288
rect -916 172968 584840 173288
rect -916 165968 584840 166288
rect -916 158968 584840 159288
rect -916 151968 584840 152288
rect -916 144968 584840 145288
rect -916 137968 584840 138288
rect -916 130968 584840 131288
rect -916 123968 584840 124288
rect -916 116968 584840 117288
rect -916 109968 584840 110288
rect -916 102968 584840 103288
rect -916 95968 584840 96288
rect -916 88968 584840 89288
rect -916 81968 584840 82288
rect -916 74968 584840 75288
rect -916 67968 584840 68288
rect -916 60968 584840 61288
rect -916 53968 584840 54288
rect -916 46968 584840 47288
rect -916 39968 584840 40288
rect -916 32968 584840 33288
rect -916 25968 584840 26288
rect -916 18968 584840 19288
rect -916 11968 584840 12288
rect -256 816 584180 1136
rect -916 156 584840 476
<< obsm5 >>
rect 12260 635608 568812 636980
rect 12260 628608 568812 634648
rect 12260 621608 568812 627648
rect 12260 614608 568812 620648
rect 12260 607608 568812 613648
rect 12260 600608 568812 606648
rect 12260 593608 568812 599648
rect 12260 586608 568812 592648
rect 12260 579608 568812 585648
rect 12260 572608 568812 578648
rect 12260 565608 568812 571648
rect 12260 558608 568812 564648
rect 12260 551608 568812 557648
rect 12260 544608 568812 550648
rect 12260 537608 568812 543648
rect 12260 530608 568812 536648
rect 12260 523608 568812 529648
rect 12260 516608 568812 522648
rect 12260 509608 568812 515648
rect 12260 502608 568812 508648
rect 12260 495608 568812 501648
rect 12260 488608 568812 494648
rect 12260 481608 568812 487648
rect 12260 474608 568812 480648
rect 12260 467608 568812 473648
rect 12260 460608 568812 466648
rect 12260 453608 568812 459648
rect 12260 446608 568812 452648
rect 12260 439608 568812 445648
rect 12260 432608 568812 438648
rect 12260 425608 568812 431648
rect 12260 418608 568812 424648
rect 12260 411608 568812 417648
rect 12260 404608 568812 410648
rect 12260 397608 568812 403648
rect 12260 390608 568812 396648
rect 12260 383608 568812 389648
rect 12260 376608 568812 382648
rect 12260 369608 568812 375648
rect 12260 362608 568812 368648
rect 12260 355608 568812 361648
rect 12260 348608 568812 354648
rect 12260 341608 568812 347648
rect 12260 334608 568812 340648
rect 12260 327608 568812 333648
rect 12260 320608 568812 326648
rect 12260 313608 568812 319648
rect 12260 306608 568812 312648
rect 12260 299608 568812 305648
rect 12260 292608 568812 298648
rect 12260 285608 568812 291648
rect 12260 278608 568812 284648
rect 12260 271608 568812 277648
rect 12260 264608 568812 270648
rect 12260 257608 568812 263648
rect 12260 250608 568812 256648
rect 12260 243608 568812 249648
rect 12260 236608 568812 242648
rect 12260 229608 568812 235648
rect 12260 222608 568812 228648
rect 12260 215608 568812 221648
rect 12260 208608 568812 214648
rect 12260 201608 568812 207648
rect 12260 194608 568812 200648
rect 12260 187608 568812 193648
rect 12260 180608 568812 186648
rect 12260 173608 568812 179648
rect 12260 166608 568812 172648
rect 12260 159608 568812 165648
rect 12260 152608 568812 158648
rect 12260 145608 568812 151648
rect 12260 138608 568812 144648
rect 12260 131608 568812 137648
rect 12260 124608 568812 130648
rect 12260 117608 568812 123648
rect 12260 110608 568812 116648
rect 12260 103608 568812 109648
rect 12260 96608 568812 102648
rect 12260 89608 568812 95648
rect 12260 82608 568812 88648
rect 12260 75608 568812 81648
rect 12260 68608 568812 74648
rect 12260 61608 568812 67648
rect 12260 54608 568812 60648
rect 12260 47608 568812 53648
rect 12260 40608 568812 46648
rect 12260 33608 568812 39648
rect 12260 26608 568812 32648
rect 12260 19608 568812 25648
rect 12260 12608 568812 18648
rect 12260 3580 568812 11648
<< labels >>
rlabel metal5 s -916 156 584840 476 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 18968 584840 19288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 32968 584840 33288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 46968 584840 47288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 60968 584840 61288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 74968 584840 75288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 88968 584840 89288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 102968 584840 103288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 116968 584840 117288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 130968 584840 131288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 144968 584840 145288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 158968 584840 159288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 172968 584840 173288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 186968 584840 187288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 200968 584840 201288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 214968 584840 215288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 228968 584840 229288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 242968 584840 243288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 256968 584840 257288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 270968 584840 271288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 284968 584840 285288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 298968 584840 299288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 312968 584840 313288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 326968 584840 327288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 340968 584840 341288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 354968 584840 355288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 368968 584840 369288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 382968 584840 383288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 396968 584840 397288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 410968 584840 411288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 424968 584840 425288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 438968 584840 439288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 452968 584840 453288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 466968 584840 467288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 480968 584840 481288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 494968 584840 495288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 508968 584840 509288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 522968 584840 523288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 536968 584840 537288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 550968 584840 551288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 564968 584840 565288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 578968 584840 579288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 592968 584840 593288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 606968 584840 607288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 620968 584840 621288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 634968 584840 635288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 648968 584840 649288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 662968 584840 663288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 676968 584840 677288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 690968 584840 691288 6 VGND
port 1 nsew ground input
rlabel metal5 s -916 703460 584840 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 26944 156 27264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 40944 156 41264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 54944 156 55264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 82944 156 83264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 96944 156 97264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 110944 156 111264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 138944 156 139264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 152944 156 153264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 166944 156 167264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 194944 156 195264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 208944 156 209264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 222944 156 223264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 250944 156 251264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 264944 156 265264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 278944 156 279264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 306944 156 307264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 320944 156 321264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 334944 156 335264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 362944 156 363264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 376944 156 377264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 390944 156 391264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 418944 156 419264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 432944 156 433264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 446944 156 447264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 474944 156 475264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 488944 156 489264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 502944 156 503264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 530944 156 531264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 544944 156 545264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 558944 156 559264 48048 6 VGND
port 1 nsew ground input
rlabel metal4 s 26944 93408 27264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 40944 93408 41264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 54944 93408 55264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 82944 93408 83264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 96944 93408 97264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 110944 93408 111264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 138944 93408 139264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 152944 93408 153264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 166944 93408 167264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 194944 93408 195264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 208944 93408 209264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 222944 93408 223264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 250944 93408 251264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 264944 93408 265264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 278944 93408 279264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 306944 93408 307264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 320944 93408 321264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 334944 93408 335264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 362944 93408 363264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 376944 93408 377264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 390944 93408 391264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 418944 93408 419264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 432944 93408 433264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 446944 93408 447264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 474944 93408 475264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 488944 93408 489264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 502944 93408 503264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 530944 93408 531264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 544944 93408 545264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 558944 93408 559264 104048 6 VGND
port 1 nsew ground input
rlabel metal4 s 26944 149408 27264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 40944 149408 41264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 54944 149408 55264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 82944 149408 83264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 96944 149408 97264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 110944 149408 111264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 138944 149408 139264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 152944 149408 153264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 166944 149408 167264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 194944 149408 195264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 208944 149408 209264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 222944 149408 223264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 250944 149408 251264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 264944 149408 265264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 278944 149408 279264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 306944 149408 307264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 320944 149408 321264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 334944 149408 335264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 362944 149408 363264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 376944 149408 377264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 390944 149408 391264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 418944 149408 419264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 432944 149408 433264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 446944 149408 447264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 474944 149408 475264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 488944 149408 489264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 502944 149408 503264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 530944 149408 531264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 544944 149408 545264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 558944 149408 559264 160048 6 VGND
port 1 nsew ground input
rlabel metal4 s 26944 205408 27264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 40944 205408 41264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 54944 205408 55264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 82944 205408 83264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 96944 205408 97264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 110944 205408 111264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 138944 205408 139264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 152944 205408 153264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 166944 205408 167264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 194944 205408 195264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 208944 205408 209264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 222944 205408 223264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 250944 205408 251264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 264944 205408 265264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 278944 205408 279264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 306944 205408 307264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 320944 205408 321264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 334944 205408 335264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 362944 205408 363264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 376944 205408 377264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 390944 205408 391264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 418944 205408 419264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 432944 205408 433264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 446944 205408 447264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 474944 205408 475264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 488944 205408 489264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 502944 205408 503264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 530944 205408 531264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 544944 205408 545264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 558944 205408 559264 216048 6 VGND
port 1 nsew ground input
rlabel metal4 s 26944 261408 27264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 40944 261408 41264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 54944 261408 55264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 82944 261408 83264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 96944 261408 97264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 110944 261408 111264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 138944 261408 139264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 152944 261408 153264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 166944 261408 167264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 194944 261408 195264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 208944 261408 209264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 222944 261408 223264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 250944 261408 251264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 264944 261408 265264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 278944 261408 279264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 306944 261408 307264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 320944 261408 321264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 334944 261408 335264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 362944 261408 363264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 376944 261408 377264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 390944 261408 391264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 418944 261408 419264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 432944 261408 433264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 446944 261408 447264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 474944 261408 475264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 488944 261408 489264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 502944 261408 503264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 530944 261408 531264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 544944 261408 545264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 558944 261408 559264 272048 6 VGND
port 1 nsew ground input
rlabel metal4 s 26944 317408 27264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 40944 317408 41264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 54944 317408 55264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 82944 317408 83264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 96944 317408 97264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 110944 317408 111264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 138944 317408 139264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 152944 317408 153264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 166944 317408 167264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 194944 317408 195264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 208944 317408 209264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 222944 317408 223264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 250944 317408 251264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 264944 317408 265264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 278944 317408 279264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 306944 317408 307264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 320944 317408 321264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 334944 317408 335264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 362944 317408 363264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 376944 317408 377264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 390944 317408 391264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 418944 317408 419264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 432944 317408 433264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 446944 317408 447264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 474944 317408 475264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 488944 317408 489264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 502944 317408 503264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 530944 317408 531264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 544944 317408 545264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 558944 317408 559264 328048 6 VGND
port 1 nsew ground input
rlabel metal4 s 26944 373408 27264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 40944 373408 41264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 54944 373408 55264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 82944 373408 83264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 96944 373408 97264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 110944 373408 111264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 138944 373408 139264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 152944 373408 153264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 166944 373408 167264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 194944 373408 195264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 208944 373408 209264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 222944 373408 223264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 250944 373408 251264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 264944 373408 265264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 278944 373408 279264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 306944 373408 307264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 320944 373408 321264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 334944 373408 335264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 362944 373408 363264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 376944 373408 377264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 390944 373408 391264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 418944 373408 419264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 432944 373408 433264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 446944 373408 447264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 474944 373408 475264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 488944 373408 489264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 502944 373408 503264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 530944 373408 531264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 544944 373408 545264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 558944 373408 559264 384048 6 VGND
port 1 nsew ground input
rlabel metal4 s 26944 429408 27264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 40944 429408 41264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 54944 429408 55264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 82944 429408 83264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 96944 429408 97264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 110944 429408 111264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 138944 429408 139264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 152944 429408 153264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 166944 429408 167264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 194944 429408 195264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 208944 429408 209264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 222944 429408 223264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 250944 429408 251264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 264944 429408 265264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 278944 429408 279264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 306944 429408 307264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 320944 429408 321264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 334944 429408 335264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 362944 429408 363264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 376944 429408 377264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 390944 429408 391264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 418944 429408 419264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 432944 429408 433264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 446944 429408 447264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 474944 429408 475264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 488944 429408 489264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 502944 429408 503264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 530944 429408 531264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 544944 429408 545264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 558944 429408 559264 440048 6 VGND
port 1 nsew ground input
rlabel metal4 s 26944 485408 27264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 40944 485408 41264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 54944 485408 55264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 82944 485408 83264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 96944 485408 97264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 110944 485408 111264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 138944 485408 139264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 152944 485408 153264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 166944 485408 167264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 194944 485408 195264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 208944 485408 209264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 222944 485408 223264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 250944 485408 251264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 264944 485408 265264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 278944 485408 279264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 306944 485408 307264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 320944 485408 321264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 334944 485408 335264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 362944 485408 363264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 376944 485408 377264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 390944 485408 391264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 418944 485408 419264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 432944 485408 433264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 446944 485408 447264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 474944 485408 475264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 488944 485408 489264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 502944 485408 503264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 530944 485408 531264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 544944 485408 545264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 558944 485408 559264 496048 6 VGND
port 1 nsew ground input
rlabel metal4 s 26944 541408 27264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 40944 541408 41264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 54944 541408 55264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 82944 541408 83264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 96944 541408 97264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 110944 541408 111264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 138944 541408 139264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 152944 541408 153264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 166944 541408 167264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 194944 541408 195264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 208944 541408 209264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 222944 541408 223264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 250944 541408 251264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 264944 541408 265264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 278944 541408 279264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 306944 541408 307264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 320944 541408 321264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 334944 541408 335264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 362944 541408 363264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 376944 541408 377264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 390944 541408 391264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 418944 541408 419264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 432944 541408 433264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 446944 541408 447264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 474944 541408 475264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 488944 541408 489264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 502944 541408 503264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 530944 541408 531264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 544944 541408 545264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 558944 541408 559264 552048 6 VGND
port 1 nsew ground input
rlabel metal4 s 26944 597408 27264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 40944 597408 41264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 54944 597408 55264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 82944 597408 83264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 96944 597408 97264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 110944 597408 111264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 138944 597408 139264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 152944 597408 153264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 166944 597408 167264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 194944 597408 195264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 208944 597408 209264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 222944 597408 223264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 250944 597408 251264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 264944 597408 265264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 278944 597408 279264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 306944 597408 307264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 320944 597408 321264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 334944 597408 335264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 362944 597408 363264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 376944 597408 377264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 390944 597408 391264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 418944 597408 419264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 432944 597408 433264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 446944 597408 447264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 474944 597408 475264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 488944 597408 489264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 502944 597408 503264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 530944 597408 531264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 544944 597408 545264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s 558944 597408 559264 608048 6 VGND
port 1 nsew ground input
rlabel metal4 s -916 156 -596 703780 4 VGND
port 1 nsew ground input
rlabel metal4 s 12944 156 13264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 26944 653408 27264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 40944 653408 41264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 54944 653408 55264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 68944 156 69264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 82944 653408 83264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 96944 653408 97264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 110944 653408 111264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 124944 156 125264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 138944 653408 139264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 152944 653408 153264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 166944 653408 167264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 180944 156 181264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 194944 653408 195264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 208944 653408 209264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 222944 653408 223264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 236944 156 237264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 250944 653408 251264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 264944 653408 265264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 278944 653408 279264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 292944 156 293264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 306944 653408 307264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 320944 653408 321264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 334944 653408 335264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 348944 156 349264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 362944 653408 363264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 376944 653408 377264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 390944 653408 391264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 404944 156 405264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 418944 653408 419264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 432944 653408 433264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 446944 653408 447264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 460944 156 461264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 474944 653408 475264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 488944 653408 489264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 502944 653408 503264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 516944 156 517264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 530944 653408 531264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 544944 653408 545264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 558944 653408 559264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 572944 156 573264 703780 6 VGND
port 1 nsew ground input
rlabel metal4 s 584520 156 584840 703780 6 VGND
port 1 nsew ground input
rlabel metal5 s -256 816 584180 1136 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 11968 584840 12288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 25968 584840 26288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 39968 584840 40288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 53968 584840 54288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 67968 584840 68288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 81968 584840 82288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 95968 584840 96288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 109968 584840 110288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 123968 584840 124288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 137968 584840 138288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 151968 584840 152288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 165968 584840 166288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 179968 584840 180288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 193968 584840 194288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 207968 584840 208288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 221968 584840 222288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 235968 584840 236288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 249968 584840 250288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 263968 584840 264288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 277968 584840 278288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 291968 584840 292288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 305968 584840 306288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 319968 584840 320288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 333968 584840 334288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 347968 584840 348288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 361968 584840 362288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 375968 584840 376288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 389968 584840 390288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 403968 584840 404288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 417968 584840 418288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 431968 584840 432288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 445968 584840 446288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 459968 584840 460288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 473968 584840 474288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 487968 584840 488288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 501968 584840 502288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 515968 584840 516288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 529968 584840 530288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 543968 584840 544288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 557968 584840 558288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 571968 584840 572288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 585968 584840 586288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 599968 584840 600288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 613968 584840 614288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 627968 584840 628288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 641968 584840 642288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 655968 584840 656288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 669968 584840 670288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 683968 584840 684288 6 VPWR
port 2 nsew power input
rlabel metal5 s -916 697968 584840 698288 6 VPWR
port 2 nsew power input
rlabel metal5 s -256 702800 584180 703120 6 VPWR
port 2 nsew power input
rlabel metal4 s 19944 156 20264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 33944 156 34264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 47944 156 48264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 75944 156 76264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 89944 156 90264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 103944 156 104264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 131944 156 132264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 145944 156 146264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 159944 156 160264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 187944 156 188264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 201944 156 202264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 215944 156 216264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 243944 156 244264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 257944 156 258264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 271944 156 272264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 299944 156 300264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 313944 156 314264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 327944 156 328264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 355944 156 356264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 369944 156 370264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 383944 156 384264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 411944 156 412264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 425944 156 426264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 439944 156 440264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 467944 156 468264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 481944 156 482264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 495944 156 496264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 523944 156 524264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 537944 156 538264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 551944 156 552264 48048 6 VPWR
port 2 nsew power input
rlabel metal4 s 19944 93408 20264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 33944 93408 34264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 47944 93408 48264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 75944 93408 76264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 89944 93408 90264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 103944 93408 104264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 131944 93408 132264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 145944 93408 146264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 159944 93408 160264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 187944 93408 188264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 201944 93408 202264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 215944 93408 216264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 243944 93408 244264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 257944 93408 258264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 271944 93408 272264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 299944 93408 300264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 313944 93408 314264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 327944 93408 328264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 355944 93408 356264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 369944 93408 370264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 383944 93408 384264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 411944 93408 412264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 425944 93408 426264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 439944 93408 440264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 467944 93408 468264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 481944 93408 482264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 495944 93408 496264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 523944 93408 524264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 537944 93408 538264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 551944 93408 552264 104048 6 VPWR
port 2 nsew power input
rlabel metal4 s 19944 149408 20264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 33944 149408 34264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 47944 149408 48264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 75944 149408 76264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 89944 149408 90264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 103944 149408 104264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 131944 149408 132264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 145944 149408 146264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 159944 149408 160264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 187944 149408 188264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 201944 149408 202264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 215944 149408 216264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 243944 149408 244264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 257944 149408 258264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 271944 149408 272264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 299944 149408 300264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 313944 149408 314264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 327944 149408 328264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 355944 149408 356264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 369944 149408 370264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 383944 149408 384264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 411944 149408 412264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 425944 149408 426264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 439944 149408 440264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 467944 149408 468264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 481944 149408 482264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 495944 149408 496264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 523944 149408 524264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 537944 149408 538264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 551944 149408 552264 160048 6 VPWR
port 2 nsew power input
rlabel metal4 s 19944 205408 20264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 33944 205408 34264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 47944 205408 48264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 75944 205408 76264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 89944 205408 90264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 103944 205408 104264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 131944 205408 132264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 145944 205408 146264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 159944 205408 160264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 187944 205408 188264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 201944 205408 202264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 215944 205408 216264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 243944 205408 244264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 257944 205408 258264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 271944 205408 272264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 299944 205408 300264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 313944 205408 314264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 327944 205408 328264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 355944 205408 356264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 369944 205408 370264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 383944 205408 384264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 411944 205408 412264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 425944 205408 426264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 439944 205408 440264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 467944 205408 468264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 481944 205408 482264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 495944 205408 496264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 523944 205408 524264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 537944 205408 538264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 551944 205408 552264 216048 6 VPWR
port 2 nsew power input
rlabel metal4 s 19944 261408 20264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 33944 261408 34264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 47944 261408 48264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 75944 261408 76264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 89944 261408 90264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 103944 261408 104264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 131944 261408 132264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 145944 261408 146264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 159944 261408 160264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 187944 261408 188264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 201944 261408 202264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 215944 261408 216264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 243944 261408 244264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 257944 261408 258264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 271944 261408 272264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 299944 261408 300264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 313944 261408 314264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 327944 261408 328264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 355944 261408 356264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 369944 261408 370264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 383944 261408 384264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 411944 261408 412264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 425944 261408 426264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 439944 261408 440264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 467944 261408 468264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 481944 261408 482264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 495944 261408 496264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 523944 261408 524264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 537944 261408 538264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 551944 261408 552264 272048 6 VPWR
port 2 nsew power input
rlabel metal4 s 19944 317408 20264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 33944 317408 34264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 47944 317408 48264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 75944 317408 76264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 89944 317408 90264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 103944 317408 104264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 131944 317408 132264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 145944 317408 146264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 159944 317408 160264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 187944 317408 188264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 201944 317408 202264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 215944 317408 216264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 243944 317408 244264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 257944 317408 258264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 271944 317408 272264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 299944 317408 300264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 313944 317408 314264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 327944 317408 328264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 355944 317408 356264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 369944 317408 370264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 383944 317408 384264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 411944 317408 412264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 425944 317408 426264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 439944 317408 440264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 467944 317408 468264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 481944 317408 482264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 495944 317408 496264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 523944 317408 524264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 537944 317408 538264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 551944 317408 552264 328048 6 VPWR
port 2 nsew power input
rlabel metal4 s 19944 373408 20264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 33944 373408 34264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 47944 373408 48264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 75944 373408 76264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 89944 373408 90264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 103944 373408 104264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 131944 373408 132264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 145944 373408 146264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 159944 373408 160264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 187944 373408 188264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 201944 373408 202264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 215944 373408 216264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 243944 373408 244264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 257944 373408 258264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 271944 373408 272264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 299944 373408 300264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 313944 373408 314264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 327944 373408 328264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 355944 373408 356264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 369944 373408 370264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 383944 373408 384264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 411944 373408 412264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 425944 373408 426264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 439944 373408 440264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 467944 373408 468264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 481944 373408 482264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 495944 373408 496264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 523944 373408 524264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 537944 373408 538264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 551944 373408 552264 384048 6 VPWR
port 2 nsew power input
rlabel metal4 s 19944 429408 20264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 33944 429408 34264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 47944 429408 48264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 75944 429408 76264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 89944 429408 90264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 103944 429408 104264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 131944 429408 132264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 145944 429408 146264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 159944 429408 160264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 187944 429408 188264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 201944 429408 202264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 215944 429408 216264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 243944 429408 244264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 257944 429408 258264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 271944 429408 272264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 299944 429408 300264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 313944 429408 314264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 327944 429408 328264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 355944 429408 356264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 369944 429408 370264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 383944 429408 384264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 411944 429408 412264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 425944 429408 426264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 439944 429408 440264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 467944 429408 468264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 481944 429408 482264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 495944 429408 496264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 523944 429408 524264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 537944 429408 538264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 551944 429408 552264 440048 6 VPWR
port 2 nsew power input
rlabel metal4 s 19944 485408 20264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 33944 485408 34264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 47944 485408 48264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 75944 485408 76264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 89944 485408 90264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 103944 485408 104264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 131944 485408 132264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 145944 485408 146264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 159944 485408 160264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 187944 485408 188264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 201944 485408 202264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 215944 485408 216264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 243944 485408 244264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 257944 485408 258264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 271944 485408 272264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 299944 485408 300264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 313944 485408 314264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 327944 485408 328264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 355944 485408 356264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 369944 485408 370264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 383944 485408 384264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 411944 485408 412264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 425944 485408 426264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 439944 485408 440264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 467944 485408 468264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 481944 485408 482264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 495944 485408 496264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 523944 485408 524264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 537944 485408 538264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 551944 485408 552264 496048 6 VPWR
port 2 nsew power input
rlabel metal4 s 19944 541408 20264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 33944 541408 34264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 47944 541408 48264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 75944 541408 76264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 89944 541408 90264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 103944 541408 104264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 131944 541408 132264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 145944 541408 146264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 159944 541408 160264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 187944 541408 188264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 201944 541408 202264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 215944 541408 216264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 243944 541408 244264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 257944 541408 258264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 271944 541408 272264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 299944 541408 300264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 313944 541408 314264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 327944 541408 328264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 355944 541408 356264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 369944 541408 370264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 383944 541408 384264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 411944 541408 412264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 425944 541408 426264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 439944 541408 440264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 467944 541408 468264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 481944 541408 482264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 495944 541408 496264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 523944 541408 524264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 537944 541408 538264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 551944 541408 552264 552048 6 VPWR
port 2 nsew power input
rlabel metal4 s 19944 597408 20264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 33944 597408 34264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 47944 597408 48264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 75944 597408 76264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 89944 597408 90264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 103944 597408 104264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 131944 597408 132264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 145944 597408 146264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 159944 597408 160264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 187944 597408 188264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 201944 597408 202264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 215944 597408 216264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 243944 597408 244264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 257944 597408 258264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 271944 597408 272264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 299944 597408 300264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 313944 597408 314264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 327944 597408 328264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 355944 597408 356264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 369944 597408 370264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 383944 597408 384264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 411944 597408 412264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 425944 597408 426264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 439944 597408 440264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 467944 597408 468264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 481944 597408 482264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 495944 597408 496264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 523944 597408 524264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 537944 597408 538264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s 551944 597408 552264 608048 6 VPWR
port 2 nsew power input
rlabel metal4 s -256 816 64 703120 4 VPWR
port 2 nsew power input
rlabel metal4 s 583860 816 584180 703120 6 VPWR
port 2 nsew power input
rlabel metal4 s 5944 156 6264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 19944 653408 20264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 33944 653408 34264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 47944 653408 48264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 61944 156 62264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 75944 653408 76264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 89944 653408 90264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 103944 653408 104264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 117944 156 118264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 131944 653408 132264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 145944 653408 146264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 159944 653408 160264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 173944 156 174264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 187944 653408 188264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 201944 653408 202264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 215944 653408 216264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 229944 156 230264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 243944 653408 244264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 257944 653408 258264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 271944 653408 272264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 285944 156 286264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 299944 653408 300264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 313944 653408 314264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 327944 653408 328264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 341944 156 342264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 355944 653408 356264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 369944 653408 370264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 383944 653408 384264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 397944 156 398264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 411944 653408 412264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 425944 653408 426264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 439944 653408 440264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 453944 156 454264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 467944 653408 468264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 481944 653408 482264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 495944 653408 496264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 509944 156 510264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 523944 653408 524264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 537944 653408 538264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 551944 653408 552264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 565944 156 566264 703780 6 VPWR
port 2 nsew power input
rlabel metal4 s 579944 156 580264 703780 6 VPWR
port 2 nsew power input
rlabel metal3 s 583200 285336 584000 285456 6 analog_io[0]
port 3 nsew signal bidirectional
rlabel metal2 s 446126 703200 446182 704000 6 analog_io[10]
port 4 nsew signal bidirectional
rlabel metal2 s 381174 703200 381230 704000 6 analog_io[11]
port 5 nsew signal bidirectional
rlabel metal2 s 316314 703200 316370 704000 6 analog_io[12]
port 6 nsew signal bidirectional
rlabel metal2 s 251454 703200 251510 704000 6 analog_io[13]
port 7 nsew signal bidirectional
rlabel metal2 s 186502 703200 186558 704000 6 analog_io[14]
port 8 nsew signal bidirectional
rlabel metal2 s 121642 703200 121698 704000 6 analog_io[15]
port 9 nsew signal bidirectional
rlabel metal2 s 56782 703200 56838 704000 6 analog_io[16]
port 10 nsew signal bidirectional
rlabel metal3 s 0 697280 800 697400 6 analog_io[17]
port 11 nsew signal bidirectional
rlabel metal3 s 0 645056 800 645176 6 analog_io[18]
port 12 nsew signal bidirectional
rlabel metal3 s 0 592968 800 593088 6 analog_io[19]
port 13 nsew signal bidirectional
rlabel metal3 s 583200 338512 584000 338632 6 analog_io[1]
port 14 nsew signal bidirectional
rlabel metal3 s 0 540744 800 540864 6 analog_io[20]
port 15 nsew signal bidirectional
rlabel metal3 s 0 488656 800 488776 6 analog_io[21]
port 16 nsew signal bidirectional
rlabel metal3 s 0 436568 800 436688 6 analog_io[22]
port 17 nsew signal bidirectional
rlabel metal3 s 0 384344 800 384464 6 analog_io[23]
port 18 nsew signal bidirectional
rlabel metal3 s 0 332256 800 332376 6 analog_io[24]
port 19 nsew signal bidirectional
rlabel metal3 s 0 280032 800 280152 6 analog_io[25]
port 20 nsew signal bidirectional
rlabel metal3 s 0 227944 800 228064 6 analog_io[26]
port 21 nsew signal bidirectional
rlabel metal3 s 0 175856 800 175976 6 analog_io[27]
port 22 nsew signal bidirectional
rlabel metal3 s 0 123632 800 123752 6 analog_io[28]
port 23 nsew signal bidirectional
rlabel metal3 s 583200 391688 584000 391808 6 analog_io[2]
port 24 nsew signal bidirectional
rlabel metal3 s 583200 444728 584000 444848 6 analog_io[3]
port 25 nsew signal bidirectional
rlabel metal3 s 583200 497904 584000 498024 6 analog_io[4]
port 26 nsew signal bidirectional
rlabel metal3 s 583200 551080 584000 551200 6 analog_io[5]
port 27 nsew signal bidirectional
rlabel metal3 s 583200 604120 584000 604240 6 analog_io[6]
port 28 nsew signal bidirectional
rlabel metal3 s 583200 657296 584000 657416 6 analog_io[7]
port 29 nsew signal bidirectional
rlabel metal2 s 575846 703200 575902 704000 6 analog_io[8]
port 30 nsew signal bidirectional
rlabel metal2 s 510986 703200 511042 704000 6 analog_io[9]
port 31 nsew signal bidirectional
rlabel metal3 s 583200 6536 584000 6656 6 io_in[0]
port 32 nsew signal input
rlabel metal3 s 583200 458056 584000 458176 6 io_in[10]
port 33 nsew signal input
rlabel metal3 s 583200 511232 584000 511352 6 io_in[11]
port 34 nsew signal input
rlabel metal3 s 583200 564272 584000 564392 6 io_in[12]
port 35 nsew signal input
rlabel metal3 s 583200 617448 584000 617568 6 io_in[13]
port 36 nsew signal input
rlabel metal3 s 583200 670624 584000 670744 6 io_in[14]
port 37 nsew signal input
rlabel metal2 s 559654 703200 559710 704000 6 io_in[15]
port 38 nsew signal input
rlabel metal2 s 494794 703200 494850 704000 6 io_in[16]
port 39 nsew signal input
rlabel metal2 s 429842 703200 429898 704000 6 io_in[17]
port 40 nsew signal input
rlabel metal2 s 364982 703200 365038 704000 6 io_in[18]
port 41 nsew signal input
rlabel metal2 s 300122 703200 300178 704000 6 io_in[19]
port 42 nsew signal input
rlabel metal3 s 583200 46248 584000 46368 6 io_in[1]
port 43 nsew signal input
rlabel metal2 s 235170 703200 235226 704000 6 io_in[20]
port 44 nsew signal input
rlabel metal2 s 170310 703200 170366 704000 6 io_in[21]
port 45 nsew signal input
rlabel metal2 s 105450 703200 105506 704000 6 io_in[22]
port 46 nsew signal input
rlabel metal2 s 40498 703200 40554 704000 6 io_in[23]
port 47 nsew signal input
rlabel metal3 s 0 684224 800 684344 6 io_in[24]
port 48 nsew signal input
rlabel metal3 s 0 632000 800 632120 6 io_in[25]
port 49 nsew signal input
rlabel metal3 s 0 579912 800 580032 6 io_in[26]
port 50 nsew signal input
rlabel metal3 s 0 527824 800 527944 6 io_in[27]
port 51 nsew signal input
rlabel metal3 s 0 475600 800 475720 6 io_in[28]
port 52 nsew signal input
rlabel metal3 s 0 423512 800 423632 6 io_in[29]
port 53 nsew signal input
rlabel metal3 s 583200 86096 584000 86216 6 io_in[2]
port 54 nsew signal input
rlabel metal3 s 0 371288 800 371408 6 io_in[30]
port 55 nsew signal input
rlabel metal3 s 0 319200 800 319320 6 io_in[31]
port 56 nsew signal input
rlabel metal3 s 0 267112 800 267232 6 io_in[32]
port 57 nsew signal input
rlabel metal3 s 0 214888 800 215008 6 io_in[33]
port 58 nsew signal input
rlabel metal3 s 0 162800 800 162920 6 io_in[34]
port 59 nsew signal input
rlabel metal3 s 0 110576 800 110696 6 io_in[35]
port 60 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 io_in[36]
port 61 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 io_in[37]
port 62 nsew signal input
rlabel metal3 s 583200 125944 584000 126064 6 io_in[3]
port 63 nsew signal input
rlabel metal3 s 583200 165792 584000 165912 6 io_in[4]
port 64 nsew signal input
rlabel metal3 s 583200 205640 584000 205760 6 io_in[5]
port 65 nsew signal input
rlabel metal3 s 583200 245488 584000 245608 6 io_in[6]
port 66 nsew signal input
rlabel metal3 s 583200 298664 584000 298784 6 io_in[7]
port 67 nsew signal input
rlabel metal3 s 583200 351840 584000 351960 6 io_in[8]
port 68 nsew signal input
rlabel metal3 s 583200 404880 584000 405000 6 io_in[9]
port 69 nsew signal input
rlabel metal3 s 583200 33056 584000 33176 6 io_oeb[0]
port 70 nsew signal output
rlabel metal3 s 583200 484576 584000 484696 6 io_oeb[10]
port 71 nsew signal output
rlabel metal3 s 583200 537752 584000 537872 6 io_oeb[11]
port 72 nsew signal output
rlabel metal3 s 583200 590928 584000 591048 6 io_oeb[12]
port 73 nsew signal output
rlabel metal3 s 583200 643968 584000 644088 6 io_oeb[13]
port 74 nsew signal output
rlabel metal3 s 583200 697144 584000 697264 6 io_oeb[14]
port 75 nsew signal output
rlabel metal2 s 527178 703200 527234 704000 6 io_oeb[15]
port 76 nsew signal output
rlabel metal2 s 462318 703200 462374 704000 6 io_oeb[16]
port 77 nsew signal output
rlabel metal2 s 397458 703200 397514 704000 6 io_oeb[17]
port 78 nsew signal output
rlabel metal2 s 332506 703200 332562 704000 6 io_oeb[18]
port 79 nsew signal output
rlabel metal2 s 267646 703200 267702 704000 6 io_oeb[19]
port 80 nsew signal output
rlabel metal3 s 583200 72904 584000 73024 6 io_oeb[1]
port 81 nsew signal output
rlabel metal2 s 202786 703200 202842 704000 6 io_oeb[20]
port 82 nsew signal output
rlabel metal2 s 137834 703200 137890 704000 6 io_oeb[21]
port 83 nsew signal output
rlabel metal2 s 72974 703200 73030 704000 6 io_oeb[22]
port 84 nsew signal output
rlabel metal2 s 8114 703200 8170 704000 6 io_oeb[23]
port 85 nsew signal output
rlabel metal3 s 0 658112 800 658232 6 io_oeb[24]
port 86 nsew signal output
rlabel metal3 s 0 606024 800 606144 6 io_oeb[25]
port 87 nsew signal output
rlabel metal3 s 0 553800 800 553920 6 io_oeb[26]
port 88 nsew signal output
rlabel metal3 s 0 501712 800 501832 6 io_oeb[27]
port 89 nsew signal output
rlabel metal3 s 0 449488 800 449608 6 io_oeb[28]
port 90 nsew signal output
rlabel metal3 s 0 397400 800 397520 6 io_oeb[29]
port 91 nsew signal output
rlabel metal3 s 583200 112752 584000 112872 6 io_oeb[2]
port 92 nsew signal output
rlabel metal3 s 0 345312 800 345432 6 io_oeb[30]
port 93 nsew signal output
rlabel metal3 s 0 293088 800 293208 6 io_oeb[31]
port 94 nsew signal output
rlabel metal3 s 0 241000 800 241120 6 io_oeb[32]
port 95 nsew signal output
rlabel metal3 s 0 188776 800 188896 6 io_oeb[33]
port 96 nsew signal output
rlabel metal3 s 0 136688 800 136808 6 io_oeb[34]
port 97 nsew signal output
rlabel metal3 s 0 84600 800 84720 6 io_oeb[35]
port 98 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 io_oeb[36]
port 99 nsew signal output
rlabel metal3 s 0 6400 800 6520 6 io_oeb[37]
port 100 nsew signal output
rlabel metal3 s 583200 152600 584000 152720 6 io_oeb[3]
port 101 nsew signal output
rlabel metal3 s 583200 192448 584000 192568 6 io_oeb[4]
port 102 nsew signal output
rlabel metal3 s 583200 232296 584000 232416 6 io_oeb[5]
port 103 nsew signal output
rlabel metal3 s 583200 272144 584000 272264 6 io_oeb[6]
port 104 nsew signal output
rlabel metal3 s 583200 325184 584000 325304 6 io_oeb[7]
port 105 nsew signal output
rlabel metal3 s 583200 378360 584000 378480 6 io_oeb[8]
port 106 nsew signal output
rlabel metal3 s 583200 431536 584000 431656 6 io_oeb[9]
port 107 nsew signal output
rlabel metal3 s 583200 19728 584000 19848 6 io_out[0]
port 108 nsew signal output
rlabel metal3 s 583200 471384 584000 471504 6 io_out[10]
port 109 nsew signal output
rlabel metal3 s 583200 524424 584000 524544 6 io_out[11]
port 110 nsew signal output
rlabel metal3 s 583200 577600 584000 577720 6 io_out[12]
port 111 nsew signal output
rlabel metal3 s 583200 630776 584000 630896 6 io_out[13]
port 112 nsew signal output
rlabel metal3 s 583200 683816 584000 683936 6 io_out[14]
port 113 nsew signal output
rlabel metal2 s 543462 703200 543518 704000 6 io_out[15]
port 114 nsew signal output
rlabel metal2 s 478510 703200 478566 704000 6 io_out[16]
port 115 nsew signal output
rlabel metal2 s 413650 703200 413706 704000 6 io_out[17]
port 116 nsew signal output
rlabel metal2 s 348790 703200 348846 704000 6 io_out[18]
port 117 nsew signal output
rlabel metal2 s 283838 703200 283894 704000 6 io_out[19]
port 118 nsew signal output
rlabel metal3 s 583200 59576 584000 59696 6 io_out[1]
port 119 nsew signal output
rlabel metal2 s 218978 703200 219034 704000 6 io_out[20]
port 120 nsew signal output
rlabel metal2 s 154118 703200 154174 704000 6 io_out[21]
port 121 nsew signal output
rlabel metal2 s 89166 703200 89222 704000 6 io_out[22]
port 122 nsew signal output
rlabel metal2 s 24306 703200 24362 704000 6 io_out[23]
port 123 nsew signal output
rlabel metal3 s 0 671168 800 671288 6 io_out[24]
port 124 nsew signal output
rlabel metal3 s 0 619080 800 619200 6 io_out[25]
port 125 nsew signal output
rlabel metal3 s 0 566856 800 566976 6 io_out[26]
port 126 nsew signal output
rlabel metal3 s 0 514768 800 514888 6 io_out[27]
port 127 nsew signal output
rlabel metal3 s 0 462544 800 462664 6 io_out[28]
port 128 nsew signal output
rlabel metal3 s 0 410456 800 410576 6 io_out[29]
port 129 nsew signal output
rlabel metal3 s 583200 99424 584000 99544 6 io_out[2]
port 130 nsew signal output
rlabel metal3 s 0 358368 800 358488 6 io_out[30]
port 131 nsew signal output
rlabel metal3 s 0 306144 800 306264 6 io_out[31]
port 132 nsew signal output
rlabel metal3 s 0 254056 800 254176 6 io_out[32]
port 133 nsew signal output
rlabel metal3 s 0 201832 800 201952 6 io_out[33]
port 134 nsew signal output
rlabel metal3 s 0 149744 800 149864 6 io_out[34]
port 135 nsew signal output
rlabel metal3 s 0 97520 800 97640 6 io_out[35]
port 136 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 io_out[36]
port 137 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 io_out[37]
port 138 nsew signal output
rlabel metal3 s 583200 139272 584000 139392 6 io_out[3]
port 139 nsew signal output
rlabel metal3 s 583200 179120 584000 179240 6 io_out[4]
port 140 nsew signal output
rlabel metal3 s 583200 218968 584000 219088 6 io_out[5]
port 141 nsew signal output
rlabel metal3 s 583200 258816 584000 258936 6 io_out[6]
port 142 nsew signal output
rlabel metal3 s 583200 311992 584000 312112 6 io_out[7]
port 143 nsew signal output
rlabel metal3 s 583200 365032 584000 365152 6 io_out[8]
port 144 nsew signal output
rlabel metal3 s 583200 418208 584000 418328 6 io_out[9]
port 145 nsew signal output
rlabel metal2 s 125874 0 125930 800 6 la_data_in[0]
port 146 nsew signal input
rlabel metal2 s 480534 0 480590 800 6 la_data_in[100]
port 147 nsew signal input
rlabel metal2 s 484030 0 484086 800 6 la_data_in[101]
port 148 nsew signal input
rlabel metal2 s 487618 0 487674 800 6 la_data_in[102]
port 149 nsew signal input
rlabel metal2 s 491114 0 491170 800 6 la_data_in[103]
port 150 nsew signal input
rlabel metal2 s 494702 0 494758 800 6 la_data_in[104]
port 151 nsew signal input
rlabel metal2 s 498198 0 498254 800 6 la_data_in[105]
port 152 nsew signal input
rlabel metal2 s 501786 0 501842 800 6 la_data_in[106]
port 153 nsew signal input
rlabel metal2 s 505374 0 505430 800 6 la_data_in[107]
port 154 nsew signal input
rlabel metal2 s 508870 0 508926 800 6 la_data_in[108]
port 155 nsew signal input
rlabel metal2 s 512458 0 512514 800 6 la_data_in[109]
port 156 nsew signal input
rlabel metal2 s 161294 0 161350 800 6 la_data_in[10]
port 157 nsew signal input
rlabel metal2 s 515954 0 516010 800 6 la_data_in[110]
port 158 nsew signal input
rlabel metal2 s 519542 0 519598 800 6 la_data_in[111]
port 159 nsew signal input
rlabel metal2 s 523038 0 523094 800 6 la_data_in[112]
port 160 nsew signal input
rlabel metal2 s 526626 0 526682 800 6 la_data_in[113]
port 161 nsew signal input
rlabel metal2 s 530122 0 530178 800 6 la_data_in[114]
port 162 nsew signal input
rlabel metal2 s 533710 0 533766 800 6 la_data_in[115]
port 163 nsew signal input
rlabel metal2 s 537206 0 537262 800 6 la_data_in[116]
port 164 nsew signal input
rlabel metal2 s 540794 0 540850 800 6 la_data_in[117]
port 165 nsew signal input
rlabel metal2 s 544382 0 544438 800 6 la_data_in[118]
port 166 nsew signal input
rlabel metal2 s 547878 0 547934 800 6 la_data_in[119]
port 167 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 la_data_in[11]
port 168 nsew signal input
rlabel metal2 s 551466 0 551522 800 6 la_data_in[120]
port 169 nsew signal input
rlabel metal2 s 554962 0 555018 800 6 la_data_in[121]
port 170 nsew signal input
rlabel metal2 s 558550 0 558606 800 6 la_data_in[122]
port 171 nsew signal input
rlabel metal2 s 562046 0 562102 800 6 la_data_in[123]
port 172 nsew signal input
rlabel metal2 s 565634 0 565690 800 6 la_data_in[124]
port 173 nsew signal input
rlabel metal2 s 569130 0 569186 800 6 la_data_in[125]
port 174 nsew signal input
rlabel metal2 s 572718 0 572774 800 6 la_data_in[126]
port 175 nsew signal input
rlabel metal2 s 576306 0 576362 800 6 la_data_in[127]
port 176 nsew signal input
rlabel metal2 s 168378 0 168434 800 6 la_data_in[12]
port 177 nsew signal input
rlabel metal2 s 171966 0 172022 800 6 la_data_in[13]
port 178 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 la_data_in[14]
port 179 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 la_data_in[15]
port 180 nsew signal input
rlabel metal2 s 182546 0 182602 800 6 la_data_in[16]
port 181 nsew signal input
rlabel metal2 s 186134 0 186190 800 6 la_data_in[17]
port 182 nsew signal input
rlabel metal2 s 189722 0 189778 800 6 la_data_in[18]
port 183 nsew signal input
rlabel metal2 s 193218 0 193274 800 6 la_data_in[19]
port 184 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 la_data_in[1]
port 185 nsew signal input
rlabel metal2 s 196806 0 196862 800 6 la_data_in[20]
port 186 nsew signal input
rlabel metal2 s 200302 0 200358 800 6 la_data_in[21]
port 187 nsew signal input
rlabel metal2 s 203890 0 203946 800 6 la_data_in[22]
port 188 nsew signal input
rlabel metal2 s 207386 0 207442 800 6 la_data_in[23]
port 189 nsew signal input
rlabel metal2 s 210974 0 211030 800 6 la_data_in[24]
port 190 nsew signal input
rlabel metal2 s 214470 0 214526 800 6 la_data_in[25]
port 191 nsew signal input
rlabel metal2 s 218058 0 218114 800 6 la_data_in[26]
port 192 nsew signal input
rlabel metal2 s 221554 0 221610 800 6 la_data_in[27]
port 193 nsew signal input
rlabel metal2 s 225142 0 225198 800 6 la_data_in[28]
port 194 nsew signal input
rlabel metal2 s 228730 0 228786 800 6 la_data_in[29]
port 195 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 la_data_in[2]
port 196 nsew signal input
rlabel metal2 s 232226 0 232282 800 6 la_data_in[30]
port 197 nsew signal input
rlabel metal2 s 235814 0 235870 800 6 la_data_in[31]
port 198 nsew signal input
rlabel metal2 s 239310 0 239366 800 6 la_data_in[32]
port 199 nsew signal input
rlabel metal2 s 242898 0 242954 800 6 la_data_in[33]
port 200 nsew signal input
rlabel metal2 s 246394 0 246450 800 6 la_data_in[34]
port 201 nsew signal input
rlabel metal2 s 249982 0 250038 800 6 la_data_in[35]
port 202 nsew signal input
rlabel metal2 s 253478 0 253534 800 6 la_data_in[36]
port 203 nsew signal input
rlabel metal2 s 257066 0 257122 800 6 la_data_in[37]
port 204 nsew signal input
rlabel metal2 s 260654 0 260710 800 6 la_data_in[38]
port 205 nsew signal input
rlabel metal2 s 264150 0 264206 800 6 la_data_in[39]
port 206 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_data_in[3]
port 207 nsew signal input
rlabel metal2 s 267738 0 267794 800 6 la_data_in[40]
port 208 nsew signal input
rlabel metal2 s 271234 0 271290 800 6 la_data_in[41]
port 209 nsew signal input
rlabel metal2 s 274822 0 274878 800 6 la_data_in[42]
port 210 nsew signal input
rlabel metal2 s 278318 0 278374 800 6 la_data_in[43]
port 211 nsew signal input
rlabel metal2 s 281906 0 281962 800 6 la_data_in[44]
port 212 nsew signal input
rlabel metal2 s 285402 0 285458 800 6 la_data_in[45]
port 213 nsew signal input
rlabel metal2 s 288990 0 289046 800 6 la_data_in[46]
port 214 nsew signal input
rlabel metal2 s 292578 0 292634 800 6 la_data_in[47]
port 215 nsew signal input
rlabel metal2 s 296074 0 296130 800 6 la_data_in[48]
port 216 nsew signal input
rlabel metal2 s 299662 0 299718 800 6 la_data_in[49]
port 217 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 la_data_in[4]
port 218 nsew signal input
rlabel metal2 s 303158 0 303214 800 6 la_data_in[50]
port 219 nsew signal input
rlabel metal2 s 306746 0 306802 800 6 la_data_in[51]
port 220 nsew signal input
rlabel metal2 s 310242 0 310298 800 6 la_data_in[52]
port 221 nsew signal input
rlabel metal2 s 313830 0 313886 800 6 la_data_in[53]
port 222 nsew signal input
rlabel metal2 s 317326 0 317382 800 6 la_data_in[54]
port 223 nsew signal input
rlabel metal2 s 320914 0 320970 800 6 la_data_in[55]
port 224 nsew signal input
rlabel metal2 s 324410 0 324466 800 6 la_data_in[56]
port 225 nsew signal input
rlabel metal2 s 327998 0 328054 800 6 la_data_in[57]
port 226 nsew signal input
rlabel metal2 s 331586 0 331642 800 6 la_data_in[58]
port 227 nsew signal input
rlabel metal2 s 335082 0 335138 800 6 la_data_in[59]
port 228 nsew signal input
rlabel metal2 s 143538 0 143594 800 6 la_data_in[5]
port 229 nsew signal input
rlabel metal2 s 338670 0 338726 800 6 la_data_in[60]
port 230 nsew signal input
rlabel metal2 s 342166 0 342222 800 6 la_data_in[61]
port 231 nsew signal input
rlabel metal2 s 345754 0 345810 800 6 la_data_in[62]
port 232 nsew signal input
rlabel metal2 s 349250 0 349306 800 6 la_data_in[63]
port 233 nsew signal input
rlabel metal2 s 352838 0 352894 800 6 la_data_in[64]
port 234 nsew signal input
rlabel metal2 s 356334 0 356390 800 6 la_data_in[65]
port 235 nsew signal input
rlabel metal2 s 359922 0 359978 800 6 la_data_in[66]
port 236 nsew signal input
rlabel metal2 s 363510 0 363566 800 6 la_data_in[67]
port 237 nsew signal input
rlabel metal2 s 367006 0 367062 800 6 la_data_in[68]
port 238 nsew signal input
rlabel metal2 s 370594 0 370650 800 6 la_data_in[69]
port 239 nsew signal input
rlabel metal2 s 147126 0 147182 800 6 la_data_in[6]
port 240 nsew signal input
rlabel metal2 s 374090 0 374146 800 6 la_data_in[70]
port 241 nsew signal input
rlabel metal2 s 377678 0 377734 800 6 la_data_in[71]
port 242 nsew signal input
rlabel metal2 s 381174 0 381230 800 6 la_data_in[72]
port 243 nsew signal input
rlabel metal2 s 384762 0 384818 800 6 la_data_in[73]
port 244 nsew signal input
rlabel metal2 s 388258 0 388314 800 6 la_data_in[74]
port 245 nsew signal input
rlabel metal2 s 391846 0 391902 800 6 la_data_in[75]
port 246 nsew signal input
rlabel metal2 s 395342 0 395398 800 6 la_data_in[76]
port 247 nsew signal input
rlabel metal2 s 398930 0 398986 800 6 la_data_in[77]
port 248 nsew signal input
rlabel metal2 s 402518 0 402574 800 6 la_data_in[78]
port 249 nsew signal input
rlabel metal2 s 406014 0 406070 800 6 la_data_in[79]
port 250 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 la_data_in[7]
port 251 nsew signal input
rlabel metal2 s 409602 0 409658 800 6 la_data_in[80]
port 252 nsew signal input
rlabel metal2 s 413098 0 413154 800 6 la_data_in[81]
port 253 nsew signal input
rlabel metal2 s 416686 0 416742 800 6 la_data_in[82]
port 254 nsew signal input
rlabel metal2 s 420182 0 420238 800 6 la_data_in[83]
port 255 nsew signal input
rlabel metal2 s 423770 0 423826 800 6 la_data_in[84]
port 256 nsew signal input
rlabel metal2 s 427266 0 427322 800 6 la_data_in[85]
port 257 nsew signal input
rlabel metal2 s 430854 0 430910 800 6 la_data_in[86]
port 258 nsew signal input
rlabel metal2 s 434442 0 434498 800 6 la_data_in[87]
port 259 nsew signal input
rlabel metal2 s 437938 0 437994 800 6 la_data_in[88]
port 260 nsew signal input
rlabel metal2 s 441526 0 441582 800 6 la_data_in[89]
port 261 nsew signal input
rlabel metal2 s 154210 0 154266 800 6 la_data_in[8]
port 262 nsew signal input
rlabel metal2 s 445022 0 445078 800 6 la_data_in[90]
port 263 nsew signal input
rlabel metal2 s 448610 0 448666 800 6 la_data_in[91]
port 264 nsew signal input
rlabel metal2 s 452106 0 452162 800 6 la_data_in[92]
port 265 nsew signal input
rlabel metal2 s 455694 0 455750 800 6 la_data_in[93]
port 266 nsew signal input
rlabel metal2 s 459190 0 459246 800 6 la_data_in[94]
port 267 nsew signal input
rlabel metal2 s 462778 0 462834 800 6 la_data_in[95]
port 268 nsew signal input
rlabel metal2 s 466274 0 466330 800 6 la_data_in[96]
port 269 nsew signal input
rlabel metal2 s 469862 0 469918 800 6 la_data_in[97]
port 270 nsew signal input
rlabel metal2 s 473450 0 473506 800 6 la_data_in[98]
port 271 nsew signal input
rlabel metal2 s 476946 0 477002 800 6 la_data_in[99]
port 272 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_data_in[9]
port 273 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_data_out[0]
port 274 nsew signal output
rlabel metal2 s 481730 0 481786 800 6 la_data_out[100]
port 275 nsew signal output
rlabel metal2 s 485226 0 485282 800 6 la_data_out[101]
port 276 nsew signal output
rlabel metal2 s 488814 0 488870 800 6 la_data_out[102]
port 277 nsew signal output
rlabel metal2 s 492310 0 492366 800 6 la_data_out[103]
port 278 nsew signal output
rlabel metal2 s 495898 0 495954 800 6 la_data_out[104]
port 279 nsew signal output
rlabel metal2 s 499394 0 499450 800 6 la_data_out[105]
port 280 nsew signal output
rlabel metal2 s 502982 0 503038 800 6 la_data_out[106]
port 281 nsew signal output
rlabel metal2 s 506478 0 506534 800 6 la_data_out[107]
port 282 nsew signal output
rlabel metal2 s 510066 0 510122 800 6 la_data_out[108]
port 283 nsew signal output
rlabel metal2 s 513562 0 513618 800 6 la_data_out[109]
port 284 nsew signal output
rlabel metal2 s 162490 0 162546 800 6 la_data_out[10]
port 285 nsew signal output
rlabel metal2 s 517150 0 517206 800 6 la_data_out[110]
port 286 nsew signal output
rlabel metal2 s 520738 0 520794 800 6 la_data_out[111]
port 287 nsew signal output
rlabel metal2 s 524234 0 524290 800 6 la_data_out[112]
port 288 nsew signal output
rlabel metal2 s 527822 0 527878 800 6 la_data_out[113]
port 289 nsew signal output
rlabel metal2 s 531318 0 531374 800 6 la_data_out[114]
port 290 nsew signal output
rlabel metal2 s 534906 0 534962 800 6 la_data_out[115]
port 291 nsew signal output
rlabel metal2 s 538402 0 538458 800 6 la_data_out[116]
port 292 nsew signal output
rlabel metal2 s 541990 0 542046 800 6 la_data_out[117]
port 293 nsew signal output
rlabel metal2 s 545486 0 545542 800 6 la_data_out[118]
port 294 nsew signal output
rlabel metal2 s 549074 0 549130 800 6 la_data_out[119]
port 295 nsew signal output
rlabel metal2 s 166078 0 166134 800 6 la_data_out[11]
port 296 nsew signal output
rlabel metal2 s 552662 0 552718 800 6 la_data_out[120]
port 297 nsew signal output
rlabel metal2 s 556158 0 556214 800 6 la_data_out[121]
port 298 nsew signal output
rlabel metal2 s 559746 0 559802 800 6 la_data_out[122]
port 299 nsew signal output
rlabel metal2 s 563242 0 563298 800 6 la_data_out[123]
port 300 nsew signal output
rlabel metal2 s 566830 0 566886 800 6 la_data_out[124]
port 301 nsew signal output
rlabel metal2 s 570326 0 570382 800 6 la_data_out[125]
port 302 nsew signal output
rlabel metal2 s 573914 0 573970 800 6 la_data_out[126]
port 303 nsew signal output
rlabel metal2 s 577410 0 577466 800 6 la_data_out[127]
port 304 nsew signal output
rlabel metal2 s 169574 0 169630 800 6 la_data_out[12]
port 305 nsew signal output
rlabel metal2 s 173162 0 173218 800 6 la_data_out[13]
port 306 nsew signal output
rlabel metal2 s 176658 0 176714 800 6 la_data_out[14]
port 307 nsew signal output
rlabel metal2 s 180246 0 180302 800 6 la_data_out[15]
port 308 nsew signal output
rlabel metal2 s 183742 0 183798 800 6 la_data_out[16]
port 309 nsew signal output
rlabel metal2 s 187330 0 187386 800 6 la_data_out[17]
port 310 nsew signal output
rlabel metal2 s 190826 0 190882 800 6 la_data_out[18]
port 311 nsew signal output
rlabel metal2 s 194414 0 194470 800 6 la_data_out[19]
port 312 nsew signal output
rlabel metal2 s 130566 0 130622 800 6 la_data_out[1]
port 313 nsew signal output
rlabel metal2 s 197910 0 197966 800 6 la_data_out[20]
port 314 nsew signal output
rlabel metal2 s 201498 0 201554 800 6 la_data_out[21]
port 315 nsew signal output
rlabel metal2 s 205086 0 205142 800 6 la_data_out[22]
port 316 nsew signal output
rlabel metal2 s 208582 0 208638 800 6 la_data_out[23]
port 317 nsew signal output
rlabel metal2 s 212170 0 212226 800 6 la_data_out[24]
port 318 nsew signal output
rlabel metal2 s 215666 0 215722 800 6 la_data_out[25]
port 319 nsew signal output
rlabel metal2 s 219254 0 219310 800 6 la_data_out[26]
port 320 nsew signal output
rlabel metal2 s 222750 0 222806 800 6 la_data_out[27]
port 321 nsew signal output
rlabel metal2 s 226338 0 226394 800 6 la_data_out[28]
port 322 nsew signal output
rlabel metal2 s 229834 0 229890 800 6 la_data_out[29]
port 323 nsew signal output
rlabel metal2 s 134154 0 134210 800 6 la_data_out[2]
port 324 nsew signal output
rlabel metal2 s 233422 0 233478 800 6 la_data_out[30]
port 325 nsew signal output
rlabel metal2 s 237010 0 237066 800 6 la_data_out[31]
port 326 nsew signal output
rlabel metal2 s 240506 0 240562 800 6 la_data_out[32]
port 327 nsew signal output
rlabel metal2 s 244094 0 244150 800 6 la_data_out[33]
port 328 nsew signal output
rlabel metal2 s 247590 0 247646 800 6 la_data_out[34]
port 329 nsew signal output
rlabel metal2 s 251178 0 251234 800 6 la_data_out[35]
port 330 nsew signal output
rlabel metal2 s 254674 0 254730 800 6 la_data_out[36]
port 331 nsew signal output
rlabel metal2 s 258262 0 258318 800 6 la_data_out[37]
port 332 nsew signal output
rlabel metal2 s 261758 0 261814 800 6 la_data_out[38]
port 333 nsew signal output
rlabel metal2 s 265346 0 265402 800 6 la_data_out[39]
port 334 nsew signal output
rlabel metal2 s 137650 0 137706 800 6 la_data_out[3]
port 335 nsew signal output
rlabel metal2 s 268842 0 268898 800 6 la_data_out[40]
port 336 nsew signal output
rlabel metal2 s 272430 0 272486 800 6 la_data_out[41]
port 337 nsew signal output
rlabel metal2 s 276018 0 276074 800 6 la_data_out[42]
port 338 nsew signal output
rlabel metal2 s 279514 0 279570 800 6 la_data_out[43]
port 339 nsew signal output
rlabel metal2 s 283102 0 283158 800 6 la_data_out[44]
port 340 nsew signal output
rlabel metal2 s 286598 0 286654 800 6 la_data_out[45]
port 341 nsew signal output
rlabel metal2 s 290186 0 290242 800 6 la_data_out[46]
port 342 nsew signal output
rlabel metal2 s 293682 0 293738 800 6 la_data_out[47]
port 343 nsew signal output
rlabel metal2 s 297270 0 297326 800 6 la_data_out[48]
port 344 nsew signal output
rlabel metal2 s 300766 0 300822 800 6 la_data_out[49]
port 345 nsew signal output
rlabel metal2 s 141238 0 141294 800 6 la_data_out[4]
port 346 nsew signal output
rlabel metal2 s 304354 0 304410 800 6 la_data_out[50]
port 347 nsew signal output
rlabel metal2 s 307942 0 307998 800 6 la_data_out[51]
port 348 nsew signal output
rlabel metal2 s 311438 0 311494 800 6 la_data_out[52]
port 349 nsew signal output
rlabel metal2 s 315026 0 315082 800 6 la_data_out[53]
port 350 nsew signal output
rlabel metal2 s 318522 0 318578 800 6 la_data_out[54]
port 351 nsew signal output
rlabel metal2 s 322110 0 322166 800 6 la_data_out[55]
port 352 nsew signal output
rlabel metal2 s 325606 0 325662 800 6 la_data_out[56]
port 353 nsew signal output
rlabel metal2 s 329194 0 329250 800 6 la_data_out[57]
port 354 nsew signal output
rlabel metal2 s 332690 0 332746 800 6 la_data_out[58]
port 355 nsew signal output
rlabel metal2 s 336278 0 336334 800 6 la_data_out[59]
port 356 nsew signal output
rlabel metal2 s 144734 0 144790 800 6 la_data_out[5]
port 357 nsew signal output
rlabel metal2 s 339866 0 339922 800 6 la_data_out[60]
port 358 nsew signal output
rlabel metal2 s 343362 0 343418 800 6 la_data_out[61]
port 359 nsew signal output
rlabel metal2 s 346950 0 347006 800 6 la_data_out[62]
port 360 nsew signal output
rlabel metal2 s 350446 0 350502 800 6 la_data_out[63]
port 361 nsew signal output
rlabel metal2 s 354034 0 354090 800 6 la_data_out[64]
port 362 nsew signal output
rlabel metal2 s 357530 0 357586 800 6 la_data_out[65]
port 363 nsew signal output
rlabel metal2 s 361118 0 361174 800 6 la_data_out[66]
port 364 nsew signal output
rlabel metal2 s 364614 0 364670 800 6 la_data_out[67]
port 365 nsew signal output
rlabel metal2 s 368202 0 368258 800 6 la_data_out[68]
port 366 nsew signal output
rlabel metal2 s 371698 0 371754 800 6 la_data_out[69]
port 367 nsew signal output
rlabel metal2 s 148322 0 148378 800 6 la_data_out[6]
port 368 nsew signal output
rlabel metal2 s 375286 0 375342 800 6 la_data_out[70]
port 369 nsew signal output
rlabel metal2 s 378874 0 378930 800 6 la_data_out[71]
port 370 nsew signal output
rlabel metal2 s 382370 0 382426 800 6 la_data_out[72]
port 371 nsew signal output
rlabel metal2 s 385958 0 386014 800 6 la_data_out[73]
port 372 nsew signal output
rlabel metal2 s 389454 0 389510 800 6 la_data_out[74]
port 373 nsew signal output
rlabel metal2 s 393042 0 393098 800 6 la_data_out[75]
port 374 nsew signal output
rlabel metal2 s 396538 0 396594 800 6 la_data_out[76]
port 375 nsew signal output
rlabel metal2 s 400126 0 400182 800 6 la_data_out[77]
port 376 nsew signal output
rlabel metal2 s 403622 0 403678 800 6 la_data_out[78]
port 377 nsew signal output
rlabel metal2 s 407210 0 407266 800 6 la_data_out[79]
port 378 nsew signal output
rlabel metal2 s 151818 0 151874 800 6 la_data_out[7]
port 379 nsew signal output
rlabel metal2 s 410798 0 410854 800 6 la_data_out[80]
port 380 nsew signal output
rlabel metal2 s 414294 0 414350 800 6 la_data_out[81]
port 381 nsew signal output
rlabel metal2 s 417882 0 417938 800 6 la_data_out[82]
port 382 nsew signal output
rlabel metal2 s 421378 0 421434 800 6 la_data_out[83]
port 383 nsew signal output
rlabel metal2 s 424966 0 425022 800 6 la_data_out[84]
port 384 nsew signal output
rlabel metal2 s 428462 0 428518 800 6 la_data_out[85]
port 385 nsew signal output
rlabel metal2 s 432050 0 432106 800 6 la_data_out[86]
port 386 nsew signal output
rlabel metal2 s 435546 0 435602 800 6 la_data_out[87]
port 387 nsew signal output
rlabel metal2 s 439134 0 439190 800 6 la_data_out[88]
port 388 nsew signal output
rlabel metal2 s 442630 0 442686 800 6 la_data_out[89]
port 389 nsew signal output
rlabel metal2 s 155406 0 155462 800 6 la_data_out[8]
port 390 nsew signal output
rlabel metal2 s 446218 0 446274 800 6 la_data_out[90]
port 391 nsew signal output
rlabel metal2 s 449806 0 449862 800 6 la_data_out[91]
port 392 nsew signal output
rlabel metal2 s 453302 0 453358 800 6 la_data_out[92]
port 393 nsew signal output
rlabel metal2 s 456890 0 456946 800 6 la_data_out[93]
port 394 nsew signal output
rlabel metal2 s 460386 0 460442 800 6 la_data_out[94]
port 395 nsew signal output
rlabel metal2 s 463974 0 464030 800 6 la_data_out[95]
port 396 nsew signal output
rlabel metal2 s 467470 0 467526 800 6 la_data_out[96]
port 397 nsew signal output
rlabel metal2 s 471058 0 471114 800 6 la_data_out[97]
port 398 nsew signal output
rlabel metal2 s 474554 0 474610 800 6 la_data_out[98]
port 399 nsew signal output
rlabel metal2 s 478142 0 478198 800 6 la_data_out[99]
port 400 nsew signal output
rlabel metal2 s 158902 0 158958 800 6 la_data_out[9]
port 401 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 la_oenb[0]
port 402 nsew signal input
rlabel metal2 s 482834 0 482890 800 6 la_oenb[100]
port 403 nsew signal input
rlabel metal2 s 486422 0 486478 800 6 la_oenb[101]
port 404 nsew signal input
rlabel metal2 s 489918 0 489974 800 6 la_oenb[102]
port 405 nsew signal input
rlabel metal2 s 493506 0 493562 800 6 la_oenb[103]
port 406 nsew signal input
rlabel metal2 s 497094 0 497150 800 6 la_oenb[104]
port 407 nsew signal input
rlabel metal2 s 500590 0 500646 800 6 la_oenb[105]
port 408 nsew signal input
rlabel metal2 s 504178 0 504234 800 6 la_oenb[106]
port 409 nsew signal input
rlabel metal2 s 507674 0 507730 800 6 la_oenb[107]
port 410 nsew signal input
rlabel metal2 s 511262 0 511318 800 6 la_oenb[108]
port 411 nsew signal input
rlabel metal2 s 514758 0 514814 800 6 la_oenb[109]
port 412 nsew signal input
rlabel metal2 s 163686 0 163742 800 6 la_oenb[10]
port 413 nsew signal input
rlabel metal2 s 518346 0 518402 800 6 la_oenb[110]
port 414 nsew signal input
rlabel metal2 s 521842 0 521898 800 6 la_oenb[111]
port 415 nsew signal input
rlabel metal2 s 525430 0 525486 800 6 la_oenb[112]
port 416 nsew signal input
rlabel metal2 s 529018 0 529074 800 6 la_oenb[113]
port 417 nsew signal input
rlabel metal2 s 532514 0 532570 800 6 la_oenb[114]
port 418 nsew signal input
rlabel metal2 s 536102 0 536158 800 6 la_oenb[115]
port 419 nsew signal input
rlabel metal2 s 539598 0 539654 800 6 la_oenb[116]
port 420 nsew signal input
rlabel metal2 s 543186 0 543242 800 6 la_oenb[117]
port 421 nsew signal input
rlabel metal2 s 546682 0 546738 800 6 la_oenb[118]
port 422 nsew signal input
rlabel metal2 s 550270 0 550326 800 6 la_oenb[119]
port 423 nsew signal input
rlabel metal2 s 167182 0 167238 800 6 la_oenb[11]
port 424 nsew signal input
rlabel metal2 s 553766 0 553822 800 6 la_oenb[120]
port 425 nsew signal input
rlabel metal2 s 557354 0 557410 800 6 la_oenb[121]
port 426 nsew signal input
rlabel metal2 s 560850 0 560906 800 6 la_oenb[122]
port 427 nsew signal input
rlabel metal2 s 564438 0 564494 800 6 la_oenb[123]
port 428 nsew signal input
rlabel metal2 s 568026 0 568082 800 6 la_oenb[124]
port 429 nsew signal input
rlabel metal2 s 571522 0 571578 800 6 la_oenb[125]
port 430 nsew signal input
rlabel metal2 s 575110 0 575166 800 6 la_oenb[126]
port 431 nsew signal input
rlabel metal2 s 578606 0 578662 800 6 la_oenb[127]
port 432 nsew signal input
rlabel metal2 s 170770 0 170826 800 6 la_oenb[12]
port 433 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_oenb[13]
port 434 nsew signal input
rlabel metal2 s 177854 0 177910 800 6 la_oenb[14]
port 435 nsew signal input
rlabel metal2 s 181442 0 181498 800 6 la_oenb[15]
port 436 nsew signal input
rlabel metal2 s 184938 0 184994 800 6 la_oenb[16]
port 437 nsew signal input
rlabel metal2 s 188526 0 188582 800 6 la_oenb[17]
port 438 nsew signal input
rlabel metal2 s 192022 0 192078 800 6 la_oenb[18]
port 439 nsew signal input
rlabel metal2 s 195610 0 195666 800 6 la_oenb[19]
port 440 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 la_oenb[1]
port 441 nsew signal input
rlabel metal2 s 199106 0 199162 800 6 la_oenb[20]
port 442 nsew signal input
rlabel metal2 s 202694 0 202750 800 6 la_oenb[21]
port 443 nsew signal input
rlabel metal2 s 206190 0 206246 800 6 la_oenb[22]
port 444 nsew signal input
rlabel metal2 s 209778 0 209834 800 6 la_oenb[23]
port 445 nsew signal input
rlabel metal2 s 213366 0 213422 800 6 la_oenb[24]
port 446 nsew signal input
rlabel metal2 s 216862 0 216918 800 6 la_oenb[25]
port 447 nsew signal input
rlabel metal2 s 220450 0 220506 800 6 la_oenb[26]
port 448 nsew signal input
rlabel metal2 s 223946 0 224002 800 6 la_oenb[27]
port 449 nsew signal input
rlabel metal2 s 227534 0 227590 800 6 la_oenb[28]
port 450 nsew signal input
rlabel metal2 s 231030 0 231086 800 6 la_oenb[29]
port 451 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 la_oenb[2]
port 452 nsew signal input
rlabel metal2 s 234618 0 234674 800 6 la_oenb[30]
port 453 nsew signal input
rlabel metal2 s 238114 0 238170 800 6 la_oenb[31]
port 454 nsew signal input
rlabel metal2 s 241702 0 241758 800 6 la_oenb[32]
port 455 nsew signal input
rlabel metal2 s 245198 0 245254 800 6 la_oenb[33]
port 456 nsew signal input
rlabel metal2 s 248786 0 248842 800 6 la_oenb[34]
port 457 nsew signal input
rlabel metal2 s 252374 0 252430 800 6 la_oenb[35]
port 458 nsew signal input
rlabel metal2 s 255870 0 255926 800 6 la_oenb[36]
port 459 nsew signal input
rlabel metal2 s 259458 0 259514 800 6 la_oenb[37]
port 460 nsew signal input
rlabel metal2 s 262954 0 263010 800 6 la_oenb[38]
port 461 nsew signal input
rlabel metal2 s 266542 0 266598 800 6 la_oenb[39]
port 462 nsew signal input
rlabel metal2 s 138846 0 138902 800 6 la_oenb[3]
port 463 nsew signal input
rlabel metal2 s 270038 0 270094 800 6 la_oenb[40]
port 464 nsew signal input
rlabel metal2 s 273626 0 273682 800 6 la_oenb[41]
port 465 nsew signal input
rlabel metal2 s 277122 0 277178 800 6 la_oenb[42]
port 466 nsew signal input
rlabel metal2 s 280710 0 280766 800 6 la_oenb[43]
port 467 nsew signal input
rlabel metal2 s 284298 0 284354 800 6 la_oenb[44]
port 468 nsew signal input
rlabel metal2 s 287794 0 287850 800 6 la_oenb[45]
port 469 nsew signal input
rlabel metal2 s 291382 0 291438 800 6 la_oenb[46]
port 470 nsew signal input
rlabel metal2 s 294878 0 294934 800 6 la_oenb[47]
port 471 nsew signal input
rlabel metal2 s 298466 0 298522 800 6 la_oenb[48]
port 472 nsew signal input
rlabel metal2 s 301962 0 302018 800 6 la_oenb[49]
port 473 nsew signal input
rlabel metal2 s 142434 0 142490 800 6 la_oenb[4]
port 474 nsew signal input
rlabel metal2 s 305550 0 305606 800 6 la_oenb[50]
port 475 nsew signal input
rlabel metal2 s 309046 0 309102 800 6 la_oenb[51]
port 476 nsew signal input
rlabel metal2 s 312634 0 312690 800 6 la_oenb[52]
port 477 nsew signal input
rlabel metal2 s 316222 0 316278 800 6 la_oenb[53]
port 478 nsew signal input
rlabel metal2 s 319718 0 319774 800 6 la_oenb[54]
port 479 nsew signal input
rlabel metal2 s 323306 0 323362 800 6 la_oenb[55]
port 480 nsew signal input
rlabel metal2 s 326802 0 326858 800 6 la_oenb[56]
port 481 nsew signal input
rlabel metal2 s 330390 0 330446 800 6 la_oenb[57]
port 482 nsew signal input
rlabel metal2 s 333886 0 333942 800 6 la_oenb[58]
port 483 nsew signal input
rlabel metal2 s 337474 0 337530 800 6 la_oenb[59]
port 484 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 la_oenb[5]
port 485 nsew signal input
rlabel metal2 s 340970 0 341026 800 6 la_oenb[60]
port 486 nsew signal input
rlabel metal2 s 344558 0 344614 800 6 la_oenb[61]
port 487 nsew signal input
rlabel metal2 s 348054 0 348110 800 6 la_oenb[62]
port 488 nsew signal input
rlabel metal2 s 351642 0 351698 800 6 la_oenb[63]
port 489 nsew signal input
rlabel metal2 s 355230 0 355286 800 6 la_oenb[64]
port 490 nsew signal input
rlabel metal2 s 358726 0 358782 800 6 la_oenb[65]
port 491 nsew signal input
rlabel metal2 s 362314 0 362370 800 6 la_oenb[66]
port 492 nsew signal input
rlabel metal2 s 365810 0 365866 800 6 la_oenb[67]
port 493 nsew signal input
rlabel metal2 s 369398 0 369454 800 6 la_oenb[68]
port 494 nsew signal input
rlabel metal2 s 372894 0 372950 800 6 la_oenb[69]
port 495 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 la_oenb[6]
port 496 nsew signal input
rlabel metal2 s 376482 0 376538 800 6 la_oenb[70]
port 497 nsew signal input
rlabel metal2 s 379978 0 380034 800 6 la_oenb[71]
port 498 nsew signal input
rlabel metal2 s 383566 0 383622 800 6 la_oenb[72]
port 499 nsew signal input
rlabel metal2 s 387154 0 387210 800 6 la_oenb[73]
port 500 nsew signal input
rlabel metal2 s 390650 0 390706 800 6 la_oenb[74]
port 501 nsew signal input
rlabel metal2 s 394238 0 394294 800 6 la_oenb[75]
port 502 nsew signal input
rlabel metal2 s 397734 0 397790 800 6 la_oenb[76]
port 503 nsew signal input
rlabel metal2 s 401322 0 401378 800 6 la_oenb[77]
port 504 nsew signal input
rlabel metal2 s 404818 0 404874 800 6 la_oenb[78]
port 505 nsew signal input
rlabel metal2 s 408406 0 408462 800 6 la_oenb[79]
port 506 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 la_oenb[7]
port 507 nsew signal input
rlabel metal2 s 411902 0 411958 800 6 la_oenb[80]
port 508 nsew signal input
rlabel metal2 s 415490 0 415546 800 6 la_oenb[81]
port 509 nsew signal input
rlabel metal2 s 418986 0 419042 800 6 la_oenb[82]
port 510 nsew signal input
rlabel metal2 s 422574 0 422630 800 6 la_oenb[83]
port 511 nsew signal input
rlabel metal2 s 426162 0 426218 800 6 la_oenb[84]
port 512 nsew signal input
rlabel metal2 s 429658 0 429714 800 6 la_oenb[85]
port 513 nsew signal input
rlabel metal2 s 433246 0 433302 800 6 la_oenb[86]
port 514 nsew signal input
rlabel metal2 s 436742 0 436798 800 6 la_oenb[87]
port 515 nsew signal input
rlabel metal2 s 440330 0 440386 800 6 la_oenb[88]
port 516 nsew signal input
rlabel metal2 s 443826 0 443882 800 6 la_oenb[89]
port 517 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_oenb[8]
port 518 nsew signal input
rlabel metal2 s 447414 0 447470 800 6 la_oenb[90]
port 519 nsew signal input
rlabel metal2 s 450910 0 450966 800 6 la_oenb[91]
port 520 nsew signal input
rlabel metal2 s 454498 0 454554 800 6 la_oenb[92]
port 521 nsew signal input
rlabel metal2 s 458086 0 458142 800 6 la_oenb[93]
port 522 nsew signal input
rlabel metal2 s 461582 0 461638 800 6 la_oenb[94]
port 523 nsew signal input
rlabel metal2 s 465170 0 465226 800 6 la_oenb[95]
port 524 nsew signal input
rlabel metal2 s 468666 0 468722 800 6 la_oenb[96]
port 525 nsew signal input
rlabel metal2 s 472254 0 472310 800 6 la_oenb[97]
port 526 nsew signal input
rlabel metal2 s 475750 0 475806 800 6 la_oenb[98]
port 527 nsew signal input
rlabel metal2 s 479338 0 479394 800 6 la_oenb[99]
port 528 nsew signal input
rlabel metal2 s 160098 0 160154 800 6 la_oenb[9]
port 529 nsew signal input
rlabel metal2 s 579802 0 579858 800 6 user_clock2
port 530 nsew signal input
rlabel metal2 s 580998 0 581054 800 6 user_irq[0]
port 531 nsew signal output
rlabel metal2 s 582194 0 582250 800 6 user_irq[1]
port 532 nsew signal output
rlabel metal2 s 583390 0 583446 800 6 user_irq[2]
port 533 nsew signal output
rlabel metal2 s 570 0 626 800 6 wb_clk_i
port 534 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wb_rst_i
port 535 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_ack_o
port 536 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 wbs_adr_i[0]
port 537 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 wbs_adr_i[10]
port 538 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 wbs_adr_i[11]
port 539 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 wbs_adr_i[12]
port 540 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 wbs_adr_i[13]
port 541 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 wbs_adr_i[14]
port 542 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 wbs_adr_i[15]
port 543 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 wbs_adr_i[16]
port 544 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 wbs_adr_i[17]
port 545 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 wbs_adr_i[18]
port 546 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 wbs_adr_i[19]
port 547 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_adr_i[1]
port 548 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 wbs_adr_i[20]
port 549 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 wbs_adr_i[21]
port 550 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 wbs_adr_i[22]
port 551 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 wbs_adr_i[23]
port 552 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 wbs_adr_i[24]
port 553 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 wbs_adr_i[25]
port 554 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 wbs_adr_i[26]
port 555 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 wbs_adr_i[27]
port 556 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 wbs_adr_i[28]
port 557 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 wbs_adr_i[29]
port 558 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_adr_i[2]
port 559 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 wbs_adr_i[30]
port 560 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 wbs_adr_i[31]
port 561 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_adr_i[3]
port 562 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 wbs_adr_i[4]
port 563 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_adr_i[5]
port 564 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_adr_i[6]
port 565 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_adr_i[7]
port 566 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 wbs_adr_i[8]
port 567 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 wbs_adr_i[9]
port 568 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_cyc_i
port 569 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_i[0]
port 570 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 wbs_dat_i[10]
port 571 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 wbs_dat_i[11]
port 572 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 wbs_dat_i[12]
port 573 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 wbs_dat_i[13]
port 574 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 wbs_dat_i[14]
port 575 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 wbs_dat_i[15]
port 576 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 wbs_dat_i[16]
port 577 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 wbs_dat_i[17]
port 578 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 wbs_dat_i[18]
port 579 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 wbs_dat_i[19]
port 580 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_i[1]
port 581 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 wbs_dat_i[20]
port 582 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 wbs_dat_i[21]
port 583 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 wbs_dat_i[22]
port 584 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 wbs_dat_i[23]
port 585 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 wbs_dat_i[24]
port 586 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 wbs_dat_i[25]
port 587 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 wbs_dat_i[26]
port 588 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 wbs_dat_i[27]
port 589 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 wbs_dat_i[28]
port 590 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 wbs_dat_i[29]
port 591 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_dat_i[2]
port 592 nsew signal input
rlabel metal2 s 119894 0 119950 800 6 wbs_dat_i[30]
port 593 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 wbs_dat_i[31]
port 594 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_i[3]
port 595 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_i[4]
port 596 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_dat_i[5]
port 597 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_dat_i[6]
port 598 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 wbs_dat_i[7]
port 599 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 wbs_dat_i[8]
port 600 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 wbs_dat_i[9]
port 601 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[0]
port 602 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 wbs_dat_o[10]
port 603 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 wbs_dat_o[11]
port 604 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 wbs_dat_o[12]
port 605 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 wbs_dat_o[13]
port 606 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 wbs_dat_o[14]
port 607 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 wbs_dat_o[15]
port 608 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 wbs_dat_o[16]
port 609 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 wbs_dat_o[17]
port 610 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 wbs_dat_o[18]
port 611 nsew signal output
rlabel metal2 s 82082 0 82138 800 6 wbs_dat_o[19]
port 612 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_o[1]
port 613 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 wbs_dat_o[20]
port 614 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 wbs_dat_o[21]
port 615 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 wbs_dat_o[22]
port 616 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 wbs_dat_o[23]
port 617 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 wbs_dat_o[24]
port 618 nsew signal output
rlabel metal2 s 103334 0 103390 800 6 wbs_dat_o[25]
port 619 nsew signal output
rlabel metal2 s 106922 0 106978 800 6 wbs_dat_o[26]
port 620 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 wbs_dat_o[27]
port 621 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 wbs_dat_o[28]
port 622 nsew signal output
rlabel metal2 s 117594 0 117650 800 6 wbs_dat_o[29]
port 623 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_o[2]
port 624 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 wbs_dat_o[30]
port 625 nsew signal output
rlabel metal2 s 124678 0 124734 800 6 wbs_dat_o[31]
port 626 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 wbs_dat_o[3]
port 627 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_o[4]
port 628 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 wbs_dat_o[5]
port 629 nsew signal output
rlabel metal2 s 35990 0 36046 800 6 wbs_dat_o[6]
port 630 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 wbs_dat_o[7]
port 631 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 wbs_dat_o[8]
port 632 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 wbs_dat_o[9]
port 633 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 wbs_sel_i[0]
port 634 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_sel_i[1]
port 635 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_sel_i[2]
port 636 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_sel_i[3]
port 637 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_stb_i
port 638 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_we_i
port 639 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 584000 704000
string LEFview TRUE
string GDS_FILE /home/egor/proj/fpga/impl/open/designs/user_project_wrapper/runs/RUN_2021.12.27_20.34.44/results/finishing/user_project_wrapper.gds
string GDS_END 442942076
string GDS_START 5213730
<< end >>

